magic
tech sky130A
magscale 1 2
timestamp 1654694770
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 348786 700544 348792 700596
rect 348844 700584 348850 700596
rect 357618 700584 357624 700596
rect 348844 700556 357624 700584
rect 348844 700544 348850 700556
rect 357618 700544 357624 700556
rect 357676 700544 357682 700596
rect 332502 700476 332508 700528
rect 332560 700516 332566 700528
rect 358906 700516 358912 700528
rect 332560 700488 358912 700516
rect 332560 700476 332566 700488
rect 358906 700476 358912 700488
rect 358964 700476 358970 700528
rect 300118 700408 300124 700460
rect 300176 700448 300182 700460
rect 357526 700448 357532 700460
rect 300176 700420 357532 700448
rect 300176 700408 300182 700420
rect 357526 700408 357532 700420
rect 357584 700408 357590 700460
rect 283834 700340 283840 700392
rect 283892 700380 283898 700392
rect 358814 700380 358820 700392
rect 283892 700352 358820 700380
rect 283892 700340 283898 700352
rect 358814 700340 358820 700352
rect 358872 700340 358878 700392
rect 105446 700272 105452 700324
rect 105504 700312 105510 700324
rect 166258 700312 166264 700324
rect 105504 700284 166264 700312
rect 105504 700272 105510 700284
rect 166258 700272 166264 700284
rect 166316 700272 166322 700324
rect 217962 700272 217968 700324
rect 218020 700312 218026 700324
rect 235166 700312 235172 700324
rect 218020 700284 235172 700312
rect 218020 700272 218026 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 357434 700312 357440 700324
rect 267700 700284 357440 700312
rect 267700 700272 267706 700284
rect 357434 700272 357440 700284
rect 357492 700272 357498 700324
rect 371878 700272 371884 700324
rect 371936 700312 371942 700324
rect 559650 700312 559656 700324
rect 371936 700284 559656 700312
rect 371936 700272 371942 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 369118 696940 369124 696992
rect 369176 696980 369182 696992
rect 580166 696980 580172 696992
rect 369176 696952 580172 696980
rect 369176 696940 369182 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 18598 670732 18604 670744
rect 3568 670704 18604 670732
rect 3568 670692 3574 670704
rect 18598 670692 18604 670704
rect 18656 670692 18662 670744
rect 360838 670692 360844 670744
rect 360896 670732 360902 670744
rect 580166 670732 580172 670744
rect 360896 670704 580172 670732
rect 360896 670692 360902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 13078 656928 13084 656940
rect 3476 656900 13084 656928
rect 3476 656888 3482 656900
rect 13078 656888 13084 656900
rect 13136 656888 13142 656940
rect 373258 643084 373264 643136
rect 373316 643124 373322 643136
rect 580166 643124 580172 643136
rect 373316 643096 580172 643124
rect 373316 643084 373322 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 197998 632108 198004 632120
rect 3476 632080 198004 632108
rect 3476 632068 3482 632080
rect 197998 632068 198004 632080
rect 198056 632068 198062 632120
rect 377398 630640 377404 630692
rect 377456 630680 377462 630692
rect 579982 630680 579988 630692
rect 377456 630652 579988 630680
rect 377456 630640 377462 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 378778 616836 378784 616888
rect 378836 616876 378842 616888
rect 580166 616876 580172 616888
rect 378836 616848 580172 616876
rect 378836 616836 378842 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 17218 605860 17224 605872
rect 3568 605832 17224 605860
rect 3568 605820 3574 605832
rect 17218 605820 17224 605832
rect 17276 605820 17282 605872
rect 363598 590656 363604 590708
rect 363656 590696 363662 590708
rect 580166 590696 580172 590708
rect 363656 590668 580172 590696
rect 363656 590656 363662 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 10318 579680 10324 579692
rect 3384 579652 10324 579680
rect 3384 579640 3390 579652
rect 10318 579640 10324 579652
rect 10376 579640 10382 579692
rect 367738 576852 367744 576904
rect 367796 576892 367802 576904
rect 580166 576892 580172 576904
rect 367796 576864 580172 576892
rect 367796 576852 367802 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 359458 563048 359464 563100
rect 359516 563088 359522 563100
rect 580166 563088 580172 563100
rect 359516 563060 580172 563088
rect 359516 563048 359522 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3142 553664 3148 553716
rect 3200 553704 3206 553716
rect 8938 553704 8944 553716
rect 3200 553676 8944 553704
rect 3200 553664 3206 553676
rect 8938 553664 8944 553676
rect 8996 553664 9002 553716
rect 500218 536800 500224 536852
rect 500276 536840 500282 536852
rect 579890 536840 579896 536852
rect 500276 536812 579896 536840
rect 500276 536800 500282 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 14458 527184 14464 527196
rect 3016 527156 14464 527184
rect 3016 527144 3022 527156
rect 14458 527144 14464 527156
rect 14516 527144 14522 527196
rect 2866 500964 2872 501016
rect 2924 501004 2930 501016
rect 21358 501004 21364 501016
rect 2924 500976 21364 501004
rect 2924 500964 2930 500976
rect 21358 500964 21364 500976
rect 21416 500964 21422 501016
rect 482278 484372 482284 484424
rect 482336 484412 482342 484424
rect 580166 484412 580172 484424
rect 482336 484384 580172 484412
rect 482336 484372 482342 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 217318 478864 217324 478916
rect 217376 478904 217382 478916
rect 220078 478904 220084 478916
rect 217376 478876 220084 478904
rect 217376 478864 217382 478876
rect 220078 478864 220084 478876
rect 220136 478864 220142 478916
rect 217594 478252 217600 478304
rect 217652 478292 217658 478304
rect 248414 478292 248420 478304
rect 217652 478264 248420 478292
rect 217652 478252 217658 478264
rect 248414 478252 248420 478264
rect 248472 478252 248478 478304
rect 309134 478252 309140 478304
rect 309192 478292 309198 478304
rect 357618 478292 357624 478304
rect 309192 478264 357624 478292
rect 309192 478252 309198 478264
rect 357618 478252 357624 478264
rect 357676 478252 357682 478304
rect 218054 478184 218060 478236
rect 218112 478224 218118 478236
rect 314746 478224 314752 478236
rect 218112 478196 314752 478224
rect 218112 478184 218118 478196
rect 314746 478184 314752 478196
rect 314804 478184 314810 478236
rect 71774 478116 71780 478168
rect 71832 478156 71838 478168
rect 346486 478156 346492 478168
rect 71832 478128 346492 478156
rect 71832 478116 71838 478128
rect 346486 478116 346492 478128
rect 346544 478116 346550 478168
rect 217502 476756 217508 476808
rect 217560 476796 217566 476808
rect 230474 476796 230480 476808
rect 217560 476768 230480 476796
rect 217560 476756 217566 476768
rect 230474 476756 230480 476768
rect 230532 476756 230538 476808
rect 238846 476756 238852 476808
rect 238904 476796 238910 476808
rect 247034 476796 247040 476808
rect 238904 476768 247040 476796
rect 238904 476756 238910 476768
rect 247034 476756 247040 476768
rect 247092 476756 247098 476808
rect 237466 476688 237472 476740
rect 237524 476728 237530 476740
rect 238754 476728 238760 476740
rect 237524 476700 238760 476728
rect 237524 476688 237530 476700
rect 238754 476688 238760 476700
rect 238812 476688 238818 476740
rect 242894 476728 242900 476740
rect 239416 476700 242900 476728
rect 233234 476620 233240 476672
rect 233292 476660 233298 476672
rect 239416 476660 239444 476700
rect 242894 476688 242900 476700
rect 242952 476688 242958 476740
rect 291194 476688 291200 476740
rect 291252 476728 291258 476740
rect 325786 476728 325792 476740
rect 291252 476700 325792 476728
rect 291252 476688 291258 476700
rect 325786 476688 325792 476700
rect 325844 476688 325850 476740
rect 249794 476660 249800 476672
rect 233292 476632 239444 476660
rect 239968 476632 249800 476660
rect 233292 476620 233298 476632
rect 233326 476552 233332 476604
rect 233384 476592 233390 476604
rect 238846 476592 238852 476604
rect 233384 476564 238852 476592
rect 233384 476552 233390 476564
rect 238846 476552 238852 476564
rect 238904 476552 238910 476604
rect 235994 476416 236000 476468
rect 236052 476456 236058 476468
rect 239968 476456 239996 476632
rect 249794 476620 249800 476632
rect 249852 476620 249858 476672
rect 251174 476620 251180 476672
rect 251232 476660 251238 476672
rect 263594 476660 263600 476672
rect 251232 476632 263600 476660
rect 251232 476620 251238 476632
rect 263594 476620 263600 476632
rect 263652 476620 263658 476672
rect 278774 476620 278780 476672
rect 278832 476660 278838 476672
rect 304994 476660 305000 476672
rect 278832 476632 305000 476660
rect 278832 476620 278838 476632
rect 304994 476620 305000 476632
rect 305052 476620 305058 476672
rect 248598 476552 248604 476604
rect 248656 476592 248662 476604
rect 260834 476592 260840 476604
rect 248656 476564 260840 476592
rect 248656 476552 248662 476564
rect 260834 476552 260840 476564
rect 260892 476552 260898 476604
rect 280154 476552 280160 476604
rect 280212 476592 280218 476604
rect 307754 476592 307760 476604
rect 280212 476564 307760 476592
rect 280212 476552 280218 476564
rect 307754 476552 307760 476564
rect 307812 476552 307818 476604
rect 242894 476484 242900 476536
rect 242952 476524 242958 476536
rect 242952 476496 244596 476524
rect 242952 476484 242958 476496
rect 236052 476428 239996 476456
rect 236052 476416 236058 476428
rect 240134 476416 240140 476468
rect 240192 476456 240198 476468
rect 240192 476428 244504 476456
rect 240192 476416 240198 476428
rect 231854 476280 231860 476332
rect 231912 476320 231918 476332
rect 235994 476320 236000 476332
rect 231912 476292 236000 476320
rect 231912 476280 231918 476292
rect 235994 476280 236000 476292
rect 236052 476280 236058 476332
rect 236086 476280 236092 476332
rect 236144 476320 236150 476332
rect 244274 476320 244280 476332
rect 236144 476292 244280 476320
rect 236144 476280 236150 476292
rect 244274 476280 244280 476292
rect 244332 476280 244338 476332
rect 238938 476212 238944 476264
rect 238996 476252 239002 476264
rect 244366 476252 244372 476264
rect 238996 476224 244372 476252
rect 238996 476212 239002 476224
rect 244366 476212 244372 476224
rect 244424 476212 244430 476264
rect 244476 476252 244504 476428
rect 244568 476388 244596 476496
rect 245746 476484 245752 476536
rect 245804 476524 245810 476536
rect 258258 476524 258264 476536
rect 245804 476496 258264 476524
rect 245804 476484 245810 476496
rect 258258 476484 258264 476496
rect 258316 476484 258322 476536
rect 259546 476484 259552 476536
rect 259604 476524 259610 476536
rect 276014 476524 276020 476536
rect 259604 476496 276020 476524
rect 259604 476484 259610 476496
rect 276014 476484 276020 476496
rect 276072 476484 276078 476536
rect 281534 476484 281540 476536
rect 281592 476524 281598 476536
rect 310514 476524 310520 476536
rect 281592 476496 310520 476524
rect 281592 476484 281598 476496
rect 310514 476484 310520 476496
rect 310572 476484 310578 476536
rect 255314 476416 255320 476468
rect 255372 476456 255378 476468
rect 268010 476456 268016 476468
rect 255372 476428 268016 476456
rect 255372 476416 255378 476428
rect 268010 476416 268016 476428
rect 268068 476416 268074 476468
rect 282914 476416 282920 476468
rect 282972 476456 282978 476468
rect 313274 476456 313280 476468
rect 282972 476428 313280 476456
rect 282972 476416 282978 476428
rect 313274 476416 313280 476428
rect 313332 476416 313338 476468
rect 244568 476360 252232 476388
rect 247310 476280 247316 476332
rect 247368 476320 247374 476332
rect 248506 476320 248512 476332
rect 247368 476292 248512 476320
rect 247368 476280 247374 476292
rect 248506 476280 248512 476292
rect 248564 476280 248570 476332
rect 252204 476320 252232 476360
rect 252554 476348 252560 476400
rect 252612 476388 252618 476400
rect 264974 476388 264980 476400
rect 252612 476360 264980 476388
rect 252612 476348 252618 476360
rect 264974 476348 264980 476360
rect 265032 476348 265038 476400
rect 284294 476348 284300 476400
rect 284352 476388 284358 476400
rect 314654 476388 314660 476400
rect 284352 476360 314660 476388
rect 284352 476348 284358 476360
rect 314654 476348 314660 476360
rect 314712 476348 314718 476400
rect 255406 476320 255412 476332
rect 252204 476292 255412 476320
rect 255406 476280 255412 476292
rect 255464 476280 255470 476332
rect 256786 476280 256792 476332
rect 256844 476320 256850 476332
rect 270494 476320 270500 476332
rect 256844 476292 270500 476320
rect 256844 476280 256850 476292
rect 270494 476280 270500 476292
rect 270552 476280 270558 476332
rect 285674 476280 285680 476332
rect 285732 476320 285738 476332
rect 317414 476320 317420 476332
rect 285732 476292 317420 476320
rect 285732 476280 285738 476292
rect 317414 476280 317420 476292
rect 317472 476280 317478 476332
rect 252738 476252 252744 476264
rect 244476 476224 252744 476252
rect 252738 476212 252744 476224
rect 252796 476212 252802 476264
rect 258166 476212 258172 476264
rect 258224 476252 258230 476264
rect 273254 476252 273260 476264
rect 258224 476224 273260 476252
rect 258224 476212 258230 476224
rect 273254 476212 273260 476224
rect 273312 476212 273318 476264
rect 288434 476212 288440 476264
rect 288492 476252 288498 476264
rect 320174 476252 320180 476264
rect 288492 476224 320180 476252
rect 288492 476212 288498 476224
rect 320174 476212 320180 476224
rect 320232 476212 320238 476264
rect 234614 476144 234620 476196
rect 234672 476184 234678 476196
rect 237374 476184 237380 476196
rect 234672 476156 237380 476184
rect 234672 476144 234678 476156
rect 237374 476144 237380 476156
rect 237432 476144 237438 476196
rect 241514 476144 241520 476196
rect 241572 476184 241578 476196
rect 245654 476184 245660 476196
rect 241572 476156 245660 476184
rect 241572 476144 241578 476156
rect 245654 476144 245660 476156
rect 245712 476144 245718 476196
rect 253842 476144 253848 476196
rect 253900 476184 253906 476196
rect 256694 476184 256700 476196
rect 253900 476156 256700 476184
rect 253900 476144 253906 476156
rect 256694 476144 256700 476156
rect 256752 476144 256758 476196
rect 260926 476144 260932 476196
rect 260984 476184 260990 476196
rect 277946 476184 277952 476196
rect 260984 476156 277952 476184
rect 260984 476144 260990 476156
rect 277946 476144 277952 476156
rect 278004 476144 278010 476196
rect 289814 476144 289820 476196
rect 289872 476184 289878 476196
rect 322934 476184 322940 476196
rect 289872 476156 322940 476184
rect 289872 476144 289878 476156
rect 322934 476144 322940 476156
rect 322992 476144 322998 476196
rect 234706 476076 234712 476128
rect 234764 476116 234770 476128
rect 235994 476116 236000 476128
rect 234764 476088 236000 476116
rect 234764 476076 234770 476088
rect 235994 476076 236000 476088
rect 236052 476076 236058 476128
rect 242802 476076 242808 476128
rect 242860 476116 242866 476128
rect 244274 476116 244280 476128
rect 242860 476088 244280 476116
rect 242860 476076 242866 476088
rect 244274 476076 244280 476088
rect 244332 476076 244338 476128
rect 245838 476076 245844 476128
rect 245896 476116 245902 476128
rect 247034 476116 247040 476128
rect 245896 476088 247040 476116
rect 245896 476076 245902 476088
rect 247034 476076 247040 476088
rect 247092 476076 247098 476128
rect 252462 476076 252468 476128
rect 252520 476116 252526 476128
rect 253934 476116 253940 476128
rect 252520 476088 253940 476116
rect 252520 476076 252526 476088
rect 253934 476076 253940 476088
rect 253992 476076 253998 476128
rect 258074 476076 258080 476128
rect 258132 476116 258138 476128
rect 262214 476116 262220 476128
rect 258132 476088 262220 476116
rect 258132 476076 258138 476088
rect 262214 476076 262220 476088
rect 262272 476076 262278 476128
rect 277578 476076 277584 476128
rect 277636 476116 277642 476128
rect 302234 476116 302240 476128
rect 277636 476088 302240 476116
rect 277636 476076 277642 476088
rect 302234 476076 302240 476088
rect 302292 476076 302298 476128
rect 219066 475328 219072 475380
rect 219124 475368 219130 475380
rect 238846 475368 238852 475380
rect 219124 475340 238852 475368
rect 219124 475328 219130 475340
rect 238846 475328 238852 475340
rect 238904 475328 238910 475380
rect 267550 475328 267556 475380
rect 267608 475368 267614 475380
rect 274634 475368 274640 475380
rect 267608 475340 274640 475368
rect 267608 475328 267614 475340
rect 274634 475328 274640 475340
rect 274692 475328 274698 475380
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 331214 474756 331220 474768
rect 3384 474728 331220 474756
rect 3384 474716 3390 474728
rect 331214 474716 331220 474728
rect 331272 474716 331278 474768
rect 219158 474036 219164 474088
rect 219216 474076 219222 474088
rect 241606 474076 241612 474088
rect 219216 474048 241612 474076
rect 219216 474036 219222 474048
rect 241606 474036 241612 474048
rect 241664 474036 241670 474088
rect 274450 474036 274456 474088
rect 274508 474076 274514 474088
rect 284386 474076 284392 474088
rect 274508 474048 284392 474076
rect 274508 474036 274514 474048
rect 284386 474036 284392 474048
rect 284444 474036 284450 474088
rect 298094 474036 298100 474088
rect 298152 474076 298158 474088
rect 377398 474076 377404 474088
rect 298152 474048 377404 474076
rect 298152 474036 298158 474048
rect 377398 474036 377404 474048
rect 377456 474036 377462 474088
rect 197998 473968 198004 474020
rect 198056 474008 198062 474020
rect 324314 474008 324320 474020
rect 198056 473980 324320 474008
rect 198056 473968 198062 473980
rect 324314 473968 324320 473980
rect 324372 473968 324378 474020
rect 217778 472676 217784 472728
rect 217836 472716 217842 472728
rect 251266 472716 251272 472728
rect 217836 472688 251272 472716
rect 217836 472676 217842 472688
rect 251266 472676 251272 472688
rect 251324 472676 251330 472728
rect 14458 472608 14464 472660
rect 14516 472648 14522 472660
rect 328454 472648 328460 472660
rect 14516 472620 328460 472648
rect 14516 472608 14522 472620
rect 328454 472608 328460 472620
rect 328512 472608 328518 472660
rect 217870 471316 217876 471368
rect 217928 471356 217934 471368
rect 254026 471356 254032 471368
rect 217928 471328 254032 471356
rect 217928 471316 217934 471328
rect 254026 471316 254032 471328
rect 254084 471316 254090 471368
rect 6914 471248 6920 471300
rect 6972 471288 6978 471300
rect 347866 471288 347872 471300
rect 6972 471260 347872 471288
rect 6972 471248 6978 471260
rect 347866 471248 347872 471260
rect 347924 471248 347930 471300
rect 300854 469888 300860 469940
rect 300912 469928 300918 469940
rect 580258 469928 580264 469940
rect 300912 469900 580264 469928
rect 300912 469888 300918 469900
rect 580258 469888 580264 469900
rect 580316 469888 580322 469940
rect 10318 469820 10324 469872
rect 10376 469860 10382 469872
rect 327074 469860 327080 469872
rect 10376 469832 327080 469860
rect 10376 469820 10382 469832
rect 327074 469820 327080 469832
rect 327132 469820 327138 469872
rect 166258 468460 166264 468512
rect 166316 468500 166322 468512
rect 317414 468500 317420 468512
rect 166316 468472 317420 468500
rect 166316 468460 166322 468472
rect 317414 468460 317420 468472
rect 317472 468460 317478 468512
rect 320174 468460 320180 468512
rect 320232 468500 320238 468512
rect 500218 468500 500224 468512
rect 320232 468472 500224 468500
rect 320232 468460 320238 468472
rect 500218 468460 500224 468472
rect 500276 468460 500282 468512
rect 295334 467168 295340 467220
rect 295392 467208 295398 467220
rect 367738 467208 367744 467220
rect 295392 467180 367744 467208
rect 295392 467168 295398 467180
rect 367738 467168 367744 467180
rect 367796 467168 367802 467220
rect 4798 467100 4804 467152
rect 4856 467140 4862 467152
rect 321554 467140 321560 467152
rect 4856 467112 321560 467140
rect 4856 467100 4862 467112
rect 321554 467100 321560 467112
rect 321612 467100 321618 467152
rect 276014 465740 276020 465792
rect 276072 465780 276078 465792
rect 300946 465780 300952 465792
rect 276072 465752 300952 465780
rect 276072 465740 276078 465752
rect 300946 465740 300952 465752
rect 301004 465740 301010 465792
rect 169754 465672 169760 465724
rect 169812 465712 169818 465724
rect 314746 465712 314752 465724
rect 169812 465684 314752 465712
rect 169812 465672 169818 465684
rect 314746 465672 314752 465684
rect 314804 465672 314810 465724
rect 318794 465672 318800 465724
rect 318852 465712 318858 465724
rect 482278 465712 482284 465724
rect 318852 465684 482284 465712
rect 318852 465672 318858 465684
rect 482278 465672 482284 465684
rect 482336 465672 482342 465724
rect 273254 464380 273260 464432
rect 273312 464420 273318 464432
rect 298186 464420 298192 464432
rect 273312 464392 298192 464420
rect 273312 464380 273318 464392
rect 298186 464380 298192 464392
rect 298244 464380 298250 464432
rect 307754 464380 307760 464432
rect 307812 464420 307818 464432
rect 364334 464420 364340 464432
rect 307812 464392 364340 464420
rect 307812 464380 307818 464392
rect 364334 464380 364340 464392
rect 364392 464380 364398 464432
rect 17218 464312 17224 464364
rect 17276 464352 17282 464364
rect 350534 464352 350540 464364
rect 17276 464324 350540 464352
rect 17276 464312 17282 464324
rect 350534 464312 350540 464324
rect 350592 464312 350598 464364
rect 266446 462952 266452 463004
rect 266504 462992 266510 463004
rect 285766 462992 285772 463004
rect 266504 462964 285772 462992
rect 266504 462952 266510 462964
rect 285766 462952 285772 462964
rect 285824 462952 285830 463004
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 332594 462380 332600 462392
rect 3384 462352 332600 462380
rect 3384 462340 3390 462352
rect 332594 462340 332600 462352
rect 332652 462340 332658 462392
rect 275922 461660 275928 461712
rect 275980 461700 275986 461712
rect 285766 461700 285772 461712
rect 275980 461672 285772 461700
rect 275980 461660 275986 461672
rect 285766 461660 285772 461672
rect 285824 461660 285830 461712
rect 219250 461592 219256 461644
rect 219308 461632 219314 461644
rect 244366 461632 244372 461644
rect 219308 461604 244372 461632
rect 219308 461592 219314 461604
rect 244366 461592 244372 461604
rect 244424 461592 244430 461644
rect 263686 461592 263692 461644
rect 263744 461632 263750 461644
rect 280246 461632 280252 461644
rect 263744 461604 280252 461632
rect 263744 461592 263750 461604
rect 280246 461592 280252 461604
rect 280304 461592 280310 461644
rect 325694 461592 325700 461644
rect 325752 461632 325758 461644
rect 373258 461632 373264 461644
rect 325752 461604 373264 461632
rect 325752 461592 325758 461604
rect 373258 461592 373264 461604
rect 373316 461592 373322 461644
rect 271874 460232 271880 460284
rect 271932 460272 271938 460284
rect 295426 460272 295432 460284
rect 271932 460244 295432 460272
rect 271932 460232 271938 460244
rect 295426 460232 295432 460244
rect 295484 460232 295490 460284
rect 322934 460232 322940 460284
rect 322992 460272 322998 460284
rect 363598 460272 363604 460284
rect 322992 460244 363604 460272
rect 322992 460232 322998 460244
rect 363598 460232 363604 460244
rect 363656 460232 363662 460284
rect 13078 460164 13084 460216
rect 13136 460204 13142 460216
rect 350626 460204 350632 460216
rect 13136 460176 350632 460204
rect 13136 460164 13142 460176
rect 350626 460164 350632 460176
rect 350684 460164 350690 460216
rect 269482 458872 269488 458924
rect 269540 458912 269546 458924
rect 289906 458912 289912 458924
rect 269540 458884 289912 458912
rect 269540 458872 269546 458884
rect 289906 458872 289912 458884
rect 289964 458872 289970 458924
rect 306374 458872 306380 458924
rect 306432 458912 306438 458924
rect 428458 458912 428464 458924
rect 306432 458884 428464 458912
rect 306432 458872 306438 458884
rect 428458 458872 428464 458884
rect 428516 458872 428522 458924
rect 8938 458804 8944 458856
rect 8996 458844 9002 458856
rect 351914 458844 351920 458856
rect 8996 458816 351920 458844
rect 8996 458804 9002 458816
rect 351914 458804 351920 458816
rect 351972 458804 351978 458856
rect 268010 457512 268016 457564
rect 268068 457552 268074 457564
rect 287054 457552 287060 457564
rect 268068 457524 287060 457552
rect 268068 457512 268074 457524
rect 287054 457512 287060 457524
rect 287112 457512 287118 457564
rect 303706 457512 303712 457564
rect 303764 457552 303770 457564
rect 494054 457552 494060 457564
rect 303764 457524 494060 457552
rect 303764 457512 303770 457524
rect 494054 457512 494060 457524
rect 494112 457512 494118 457564
rect 21358 457444 21364 457496
rect 21416 457484 21422 457496
rect 352466 457484 352472 457496
rect 21416 457456 352472 457484
rect 21416 457444 21422 457456
rect 352466 457444 352472 457456
rect 352524 457444 352530 457496
rect 265066 456084 265072 456136
rect 265124 456124 265130 456136
rect 283006 456124 283012 456136
rect 265124 456096 283012 456124
rect 265124 456084 265130 456096
rect 283006 456084 283012 456096
rect 283064 456084 283070 456136
rect 301314 456084 301320 456136
rect 301372 456124 301378 456136
rect 371878 456124 371884 456136
rect 301372 456096 371884 456124
rect 301372 456084 301378 456096
rect 371878 456084 371884 456096
rect 371936 456084 371942 456136
rect 18598 456016 18604 456068
rect 18656 456056 18662 456068
rect 323762 456056 323768 456068
rect 18656 456028 323768 456056
rect 18656 456016 18662 456028
rect 323762 456016 323768 456028
rect 323820 456016 323826 456068
rect 269022 455336 269028 455388
rect 269080 455376 269086 455388
rect 276474 455376 276480 455388
rect 269080 455348 276480 455376
rect 269080 455336 269086 455348
rect 276474 455336 276480 455348
rect 276532 455336 276538 455388
rect 274542 454724 274548 454776
rect 274600 454764 274606 454776
rect 283006 454764 283012 454776
rect 274600 454736 283012 454764
rect 274600 454724 274606 454736
rect 283006 454724 283012 454736
rect 283064 454724 283070 454776
rect 219342 454656 219348 454708
rect 219400 454696 219406 454708
rect 247126 454696 247132 454708
rect 219400 454668 247132 454696
rect 219400 454656 219406 454668
rect 247126 454656 247132 454668
rect 247184 454656 247190 454708
rect 280062 454656 280068 454708
rect 280120 454696 280126 454708
rect 290458 454696 290464 454708
rect 280120 454668 290464 454696
rect 280120 454656 280126 454668
rect 290458 454656 290464 454668
rect 290516 454656 290522 454708
rect 298922 454656 298928 454708
rect 298980 454696 298986 454708
rect 360838 454696 360844 454708
rect 298980 454668 360844 454696
rect 298980 454656 298986 454668
rect 360838 454656 360844 454668
rect 360896 454656 360902 454708
rect 267642 453364 267648 453416
rect 267700 453404 267706 453416
rect 273346 453404 273352 453416
rect 267700 453376 273352 453404
rect 267700 453364 267706 453376
rect 273346 453364 273352 453376
rect 273404 453364 273410 453416
rect 277302 453364 277308 453416
rect 277360 453404 277366 453416
rect 287330 453404 287336 453416
rect 277360 453376 287336 453404
rect 277360 453364 277366 453376
rect 287330 453364 287336 453376
rect 287388 453364 287394 453416
rect 270954 453296 270960 453348
rect 271012 453336 271018 453348
rect 292574 453336 292580 453348
rect 271012 453308 292580 453336
rect 271012 453296 271018 453308
rect 292574 453296 292580 453308
rect 292632 453296 292638 453348
rect 296714 453296 296720 453348
rect 296772 453336 296778 453348
rect 378778 453336 378784 453348
rect 296772 453308 378784 453336
rect 296772 453296 296778 453308
rect 378778 453296 378784 453308
rect 378836 453296 378842 453348
rect 271782 452752 271788 452804
rect 271840 452792 271846 452804
rect 279602 452792 279608 452804
rect 271840 452764 279608 452792
rect 271840 452752 271846 452764
rect 279602 452752 279608 452764
rect 279660 452752 279666 452804
rect 266262 451936 266268 451988
rect 266320 451976 266326 451988
rect 271966 451976 271972 451988
rect 266320 451948 271972 451976
rect 266320 451936 266326 451948
rect 271966 451936 271972 451948
rect 272024 451936 272030 451988
rect 273162 451936 273168 451988
rect 273220 451976 273226 451988
rect 281718 451976 281724 451988
rect 273220 451948 281724 451976
rect 273220 451936 273226 451948
rect 281718 451936 281724 451948
rect 281776 451936 281782 451988
rect 217686 451868 217692 451920
rect 217744 451908 217750 451920
rect 231946 451908 231952 451920
rect 217744 451880 231952 451908
rect 217744 451868 217750 451880
rect 231946 451868 231952 451880
rect 232004 451868 232010 451920
rect 270402 451868 270408 451920
rect 270460 451908 270466 451920
rect 277486 451908 277492 451920
rect 270460 451880 277492 451908
rect 270460 451868 270466 451880
rect 277486 451868 277492 451880
rect 277544 451868 277550 451920
rect 278682 451868 278688 451920
rect 278740 451908 278746 451920
rect 288802 451908 288808 451920
rect 278740 451880 288808 451908
rect 278740 451868 278746 451880
rect 288802 451868 288808 451880
rect 288860 451868 288866 451920
rect 294322 451868 294328 451920
rect 294380 451908 294386 451920
rect 359458 451908 359464 451920
rect 294380 451880 359464 451908
rect 294380 451868 294386 451880
rect 359458 451868 359464 451880
rect 359516 451868 359522 451920
rect 328086 450644 328092 450696
rect 328144 450684 328150 450696
rect 369118 450684 369124 450696
rect 328144 450656 369124 450684
rect 328144 450644 328150 450656
rect 369118 450644 369124 450656
rect 369176 450644 369182 450696
rect 3510 450576 3516 450628
rect 3568 450616 3574 450628
rect 328822 450616 328828 450628
rect 3568 450588 328828 450616
rect 3568 450576 3574 450588
rect 328822 450576 328828 450588
rect 328880 450576 328886 450628
rect 3602 450508 3608 450560
rect 3660 450548 3666 450560
rect 331214 450548 331220 450560
rect 3660 450520 331220 450548
rect 3660 450508 3666 450520
rect 331214 450508 331220 450520
rect 331272 450508 331278 450560
rect 307938 449556 307944 449608
rect 307996 449596 308002 449608
rect 412634 449596 412640 449608
rect 307996 449568 412640 449596
rect 307996 449556 308002 449568
rect 412634 449556 412640 449568
rect 412692 449556 412698 449608
rect 153194 449488 153200 449540
rect 153252 449528 153258 449540
rect 317230 449528 317236 449540
rect 153252 449500 317236 449528
rect 153252 449488 153258 449500
rect 317230 449488 317236 449500
rect 317288 449488 317294 449540
rect 305546 449420 305552 449472
rect 305604 449460 305610 449472
rect 477494 449460 477500 449472
rect 305604 449432 477500 449460
rect 305604 449420 305610 449432
rect 477494 449420 477500 449432
rect 477552 449420 477558 449472
rect 88334 449352 88340 449404
rect 88392 449392 88398 449404
rect 319530 449392 319536 449404
rect 88392 449364 319536 449392
rect 88392 449352 88398 449364
rect 319530 449352 319536 449364
rect 319588 449352 319594 449404
rect 303246 449284 303252 449336
rect 303304 449324 303310 449336
rect 542354 449324 542360 449336
rect 303304 449296 542360 449324
rect 303304 449284 303310 449296
rect 542354 449284 542360 449296
rect 542412 449284 542418 449336
rect 23474 449216 23480 449268
rect 23532 449256 23538 449268
rect 321830 449256 321836 449268
rect 23532 449228 321836 449256
rect 23532 449216 23538 449228
rect 321830 449216 321836 449228
rect 321888 449216 321894 449268
rect 3418 449148 3424 449200
rect 3476 449188 3482 449200
rect 326522 449188 326528 449200
rect 3476 449160 326528 449188
rect 3476 449148 3482 449160
rect 326522 449148 326528 449160
rect 326580 449148 326586 449200
rect 335078 448128 335084 448180
rect 335136 448168 335142 448180
rect 397454 448168 397460 448180
rect 335136 448140 397460 448168
rect 335136 448128 335142 448140
rect 397454 448128 397460 448140
rect 397512 448128 397518 448180
rect 332778 448060 332784 448112
rect 332836 448100 332842 448112
rect 462314 448100 462320 448112
rect 332836 448072 462320 448100
rect 332836 448060 332842 448072
rect 462314 448060 462320 448072
rect 462372 448060 462378 448112
rect 201494 447992 201500 448044
rect 201552 448032 201558 448044
rect 342070 448032 342076 448044
rect 201552 448004 342076 448032
rect 201552 447992 201558 448004
rect 342070 447992 342076 448004
rect 342128 447992 342134 448044
rect 136634 447924 136640 447976
rect 136692 447964 136698 447976
rect 344370 447964 344376 447976
rect 136692 447936 344376 447964
rect 136692 447924 136698 447936
rect 344370 447924 344376 447936
rect 344428 447924 344434 447976
rect 40034 447856 40040 447908
rect 40092 447896 40098 447908
rect 320358 447896 320364 447908
rect 40092 447868 320364 447896
rect 40092 447856 40098 447868
rect 320358 447856 320364 447868
rect 320416 447856 320422 447908
rect 330386 447856 330392 447908
rect 330444 447896 330450 447908
rect 527174 447896 527180 447908
rect 330444 447868 527180 447896
rect 330444 447856 330450 447868
rect 527174 447856 527180 447868
rect 527232 447856 527238 447908
rect 2866 447788 2872 447840
rect 2924 447828 2930 447840
rect 353662 447828 353668 447840
rect 2924 447800 353668 447828
rect 2924 447788 2930 447800
rect 353662 447788 353668 447800
rect 353720 447788 353726 447840
rect 231854 447040 231860 447092
rect 231912 447080 231918 447092
rect 232406 447080 232412 447092
rect 231912 447052 232412 447080
rect 231912 447040 231918 447052
rect 232406 447040 232412 447052
rect 232464 447040 232470 447092
rect 235994 447040 236000 447092
rect 236052 447080 236058 447092
rect 237006 447080 237012 447092
rect 236052 447052 237012 447080
rect 236052 447040 236058 447052
rect 237006 447040 237012 447052
rect 237064 447040 237070 447092
rect 241514 447040 241520 447092
rect 241572 447080 241578 447092
rect 242342 447080 242348 447092
rect 241572 447052 242348 447080
rect 241572 447040 241578 447052
rect 242342 447040 242348 447052
rect 242400 447040 242406 447092
rect 245746 447040 245752 447092
rect 245804 447080 245810 447092
rect 246390 447080 246396 447092
rect 245804 447052 246396 447080
rect 245804 447040 245810 447052
rect 246390 447040 246396 447052
rect 246448 447040 246454 447092
rect 248414 447040 248420 447092
rect 248472 447080 248478 447092
rect 249334 447080 249340 447092
rect 248472 447052 249340 447080
rect 248472 447040 248478 447052
rect 249334 447040 249340 447052
rect 249392 447040 249398 447092
rect 252554 447040 252560 447092
rect 252612 447080 252618 447092
rect 253198 447080 253204 447092
rect 252612 447052 253204 447080
rect 252612 447040 252618 447052
rect 253198 447040 253204 447052
rect 253256 447040 253262 447092
rect 255958 447040 255964 447092
rect 256016 447080 256022 447092
rect 258258 447080 258264 447092
rect 256016 447052 258264 447080
rect 256016 447040 256022 447052
rect 258258 447040 258264 447052
rect 258316 447040 258322 447092
rect 258718 447040 258724 447092
rect 258776 447080 258782 447092
rect 261110 447080 261116 447092
rect 258776 447052 261116 447080
rect 258776 447040 258782 447052
rect 261110 447040 261116 447052
rect 261168 447040 261174 447092
rect 262858 447040 262864 447092
rect 262916 447080 262922 447092
rect 267550 447080 267556 447092
rect 262916 447052 267556 447080
rect 262916 447040 262922 447052
rect 267550 447040 267556 447052
rect 267608 447040 267614 447092
rect 271874 447040 271880 447092
rect 271932 447080 271938 447092
rect 272702 447080 272708 447092
rect 271932 447052 272708 447080
rect 271932 447040 271938 447052
rect 272702 447040 272708 447052
rect 272760 447040 272766 447092
rect 273254 447040 273260 447092
rect 273312 447080 273318 447092
rect 274174 447080 274180 447092
rect 273312 447052 274180 447080
rect 273312 447040 273318 447052
rect 274174 447040 274180 447052
rect 274232 447040 274238 447092
rect 277486 447040 277492 447092
rect 277544 447080 277550 447092
rect 278038 447080 278044 447092
rect 277544 447052 278044 447080
rect 277544 447040 277550 447052
rect 278038 447040 278044 447052
rect 278096 447040 278102 447092
rect 281534 447040 281540 447092
rect 281592 447080 281598 447092
rect 281902 447080 281908 447092
rect 281592 447052 281908 447080
rect 281592 447040 281598 447052
rect 281902 447040 281908 447052
rect 281960 447040 281966 447092
rect 282914 447040 282920 447092
rect 282972 447080 282978 447092
rect 283558 447080 283564 447092
rect 282972 447052 283564 447080
rect 282972 447040 282978 447052
rect 283558 447040 283564 447052
rect 283616 447040 283622 447092
rect 284294 447040 284300 447092
rect 284352 447080 284358 447092
rect 285030 447080 285036 447092
rect 284352 447052 285036 447080
rect 284352 447040 284358 447052
rect 285030 447040 285036 447052
rect 285088 447040 285094 447092
rect 285674 447040 285680 447092
rect 285732 447080 285738 447092
rect 286686 447080 286692 447092
rect 285732 447052 286692 447080
rect 285732 447040 285738 447052
rect 286686 447040 286692 447052
rect 286744 447040 286750 447092
rect 350534 447040 350540 447092
rect 350592 447080 350598 447092
rect 351086 447080 351092 447092
rect 350592 447052 351092 447080
rect 350592 447040 350598 447052
rect 351086 447040 351092 447052
rect 351144 447040 351150 447092
rect 256602 446972 256608 447024
rect 256660 447012 256666 447024
rect 259822 447012 259828 447024
rect 256660 446984 259828 447012
rect 256660 446972 256666 446984
rect 259822 446972 259828 446984
rect 259880 446972 259886 447024
rect 260742 446972 260748 447024
rect 260800 447012 260806 447024
rect 264514 447012 264520 447024
rect 260800 446984 264520 447012
rect 260800 446972 260806 446984
rect 264514 446972 264520 446984
rect 264572 446972 264578 447024
rect 264238 446904 264244 446956
rect 264296 446944 264302 446956
rect 269114 446944 269120 446956
rect 264296 446916 269120 446944
rect 264296 446904 264302 446916
rect 269114 446904 269120 446916
rect 269172 446904 269178 446956
rect 57238 446768 57244 446820
rect 57296 446808 57302 446820
rect 349798 446808 349804 446820
rect 57296 446780 349804 446808
rect 57296 446768 57302 446780
rect 349798 446768 349804 446780
rect 349856 446768 349862 446820
rect 339678 446700 339684 446752
rect 339736 446740 339742 446752
rect 357434 446740 357440 446752
rect 339736 446712 357440 446740
rect 339736 446700 339742 446712
rect 357434 446700 357440 446712
rect 357492 446700 357498 446752
rect 217962 446632 217968 446684
rect 218020 446672 218026 446684
rect 313366 446672 313372 446684
rect 218020 446644 313372 446672
rect 218020 446632 218026 446644
rect 313366 446632 313372 446644
rect 313424 446632 313430 446684
rect 337378 446632 337384 446684
rect 337436 446672 337442 446684
rect 358906 446672 358912 446684
rect 337436 446644 358912 446672
rect 337436 446632 337442 446644
rect 358906 446632 358912 446644
rect 358964 446632 358970 446684
rect 312538 446564 312544 446616
rect 312596 446604 312602 446616
rect 358814 446604 358820 446616
rect 312596 446576 358820 446604
rect 312596 446564 312602 446576
rect 358814 446564 358820 446576
rect 358872 446564 358878 446616
rect 261478 446496 261484 446548
rect 261536 446536 261542 446548
rect 265986 446536 265992 446548
rect 261536 446508 265992 446536
rect 261536 446496 261542 446508
rect 265986 446496 265992 446508
rect 266044 446496 266050 446548
rect 310974 446496 310980 446548
rect 311032 446536 311038 446548
rect 357526 446536 357532 446548
rect 311032 446508 357532 446536
rect 311032 446496 311038 446508
rect 357526 446496 357532 446508
rect 357584 446496 357590 446548
rect 220078 446428 220084 446480
rect 220136 446468 220142 446480
rect 230382 446468 230388 446480
rect 220136 446440 230388 446468
rect 220136 446428 220142 446440
rect 230382 446428 230388 446440
rect 230440 446428 230446 446480
rect 265618 446428 265624 446480
rect 265676 446468 265682 446480
rect 270678 446468 270684 446480
rect 265676 446440 270684 446468
rect 265676 446428 265682 446440
rect 270678 446428 270684 446440
rect 270736 446428 270742 446480
rect 307110 446428 307116 446480
rect 307168 446468 307174 446480
rect 364978 446468 364984 446480
rect 307168 446440 364984 446468
rect 307168 446428 307174 446440
rect 364978 446428 364984 446440
rect 365036 446428 365042 446480
rect 311802 446360 311808 446412
rect 311860 446400 311866 446412
rect 362218 446400 362224 446412
rect 311860 446372 362224 446400
rect 311860 446360 311866 446372
rect 362218 446360 362224 446372
rect 362276 446360 362282 446412
rect 304810 446292 304816 446344
rect 304868 446332 304874 446344
rect 363598 446332 363604 446344
rect 304868 446304 363604 446332
rect 304868 446292 304874 446304
rect 363598 446292 363604 446304
rect 363656 446292 363662 446344
rect 293126 446224 293132 446276
rect 293184 446264 293190 446276
rect 362310 446264 362316 446276
rect 293184 446236 362316 446264
rect 293184 446224 293190 446236
rect 362310 446224 362316 446236
rect 362368 446224 362374 446276
rect 292390 446156 292396 446208
rect 292448 446196 292454 446208
rect 373258 446196 373264 446208
rect 292448 446168 373264 446196
rect 292448 446156 292454 446168
rect 373258 446156 373264 446168
rect 373316 446156 373322 446208
rect 244366 446088 244372 446140
rect 244424 446128 244430 446140
rect 345106 446128 345112 446140
rect 244424 446100 345112 446128
rect 244424 446088 244430 446100
rect 345106 446088 345112 446100
rect 345164 446088 345170 446140
rect 229830 446020 229836 446072
rect 229888 446060 229894 446072
rect 338206 446060 338212 446072
rect 229888 446032 338212 446060
rect 229888 446020 229894 446032
rect 338206 446020 338212 446032
rect 338264 446020 338270 446072
rect 228358 445952 228364 446004
rect 228416 445992 228422 446004
rect 347498 445992 347504 446004
rect 228416 445964 347504 445992
rect 228416 445952 228422 445964
rect 347498 445952 347504 445964
rect 347556 445952 347562 446004
rect 229738 445884 229744 445936
rect 229796 445924 229802 445936
rect 359918 445924 359924 445936
rect 229796 445896 359924 445924
rect 229796 445884 229802 445896
rect 359918 445884 359924 445896
rect 359976 445884 359982 445936
rect 293954 445816 293960 445868
rect 294012 445856 294018 445868
rect 458818 445856 458824 445868
rect 294012 445828 458824 445856
rect 294012 445816 294018 445828
rect 458818 445816 458824 445828
rect 458876 445816 458882 445868
rect 302510 445748 302516 445800
rect 302568 445788 302574 445800
rect 311158 445788 311164 445800
rect 302568 445760 311164 445788
rect 302568 445748 302574 445760
rect 311158 445748 311164 445760
rect 311216 445748 311222 445800
rect 316402 445748 316408 445800
rect 316460 445788 316466 445800
rect 333974 445788 333980 445800
rect 316460 445760 333980 445788
rect 316460 445748 316466 445760
rect 333974 445748 333980 445760
rect 334032 445748 334038 445800
rect 253934 445408 253940 445460
rect 253992 445448 253998 445460
rect 254854 445448 254860 445460
rect 253992 445420 254860 445448
rect 253992 445408 253998 445420
rect 254854 445408 254860 445420
rect 254912 445408 254918 445460
rect 228542 445204 228548 445256
rect 228600 445244 228606 445256
rect 336642 445244 336648 445256
rect 228600 445216 336648 445244
rect 228600 445204 228606 445216
rect 336642 445204 336648 445216
rect 336700 445204 336706 445256
rect 225690 445136 225696 445188
rect 225748 445176 225754 445188
rect 338942 445176 338948 445188
rect 225748 445148 338948 445176
rect 225748 445136 225754 445148
rect 338942 445136 338948 445148
rect 339000 445136 339006 445188
rect 333974 445068 333980 445120
rect 334032 445108 334038 445120
rect 580350 445108 580356 445120
rect 334032 445080 580356 445108
rect 334032 445068 334038 445080
rect 580350 445068 580356 445080
rect 580408 445068 580414 445120
rect 311158 445000 311164 445052
rect 311216 445040 311222 445052
rect 580258 445040 580264 445052
rect 311216 445012 580264 445040
rect 311216 445000 311222 445012
rect 580258 445000 580264 445012
rect 580316 445000 580322 445052
rect 224218 444932 224224 444984
rect 224276 444972 224282 444984
rect 341242 444972 341248 444984
rect 224276 444944 341248 444972
rect 224276 444932 224282 444944
rect 341242 444932 341248 444944
rect 341300 444932 341306 444984
rect 228450 444864 228456 444916
rect 228508 444904 228514 444916
rect 355962 444904 355968 444916
rect 228508 444876 355968 444904
rect 228508 444864 228514 444876
rect 355962 444864 355968 444876
rect 356020 444864 356026 444916
rect 300118 444796 300124 444848
rect 300176 444836 300182 444848
rect 460198 444836 460204 444848
rect 300176 444808 460204 444836
rect 300176 444796 300182 444808
rect 460198 444796 460204 444808
rect 460256 444796 460262 444848
rect 295518 444728 295524 444780
rect 295576 444768 295582 444780
rect 494698 444768 494704 444780
rect 295576 444740 494704 444768
rect 295576 444728 295582 444740
rect 494698 444728 494704 444740
rect 494756 444728 494762 444780
rect 86218 444660 86224 444712
rect 86276 444700 86282 444712
rect 343634 444700 343640 444712
rect 86276 444672 343640 444700
rect 86276 444660 86282 444672
rect 343634 444660 343640 444672
rect 343692 444660 343698 444712
rect 84838 444592 84844 444644
rect 84896 444632 84902 444644
rect 345934 444632 345940 444644
rect 84896 444604 345940 444632
rect 84896 444592 84902 444604
rect 345934 444592 345940 444604
rect 345992 444592 345998 444644
rect 82078 444524 82084 444576
rect 82136 444564 82142 444576
rect 348234 444564 348240 444576
rect 82136 444536 348240 444564
rect 82136 444524 82142 444536
rect 348234 444524 348240 444536
rect 348292 444524 348298 444576
rect 80698 444456 80704 444508
rect 80756 444496 80762 444508
rect 358354 444496 358360 444508
rect 80756 444468 358360 444496
rect 80756 444456 80762 444468
rect 358354 444456 358360 444468
rect 358412 444456 358418 444508
rect 7558 444388 7564 444440
rect 7616 444428 7622 444440
rect 334250 444428 334256 444440
rect 7616 444400 334256 444428
rect 7616 444388 7622 444400
rect 334250 444388 334256 444400
rect 334308 444388 334314 444440
rect 309502 443708 309508 443760
rect 309560 443748 309566 443760
rect 309560 443720 311894 443748
rect 309560 443708 309566 443720
rect 3510 443640 3516 443692
rect 3568 443680 3574 443692
rect 244366 443680 244372 443692
rect 3568 443652 244372 443680
rect 3568 443640 3574 443652
rect 244366 443640 244372 443652
rect 244424 443640 244430 443692
rect 311866 443612 311894 443720
rect 314378 443640 314384 443692
rect 314436 443680 314442 443692
rect 369118 443680 369124 443692
rect 314436 443652 369124 443680
rect 314436 443640 314442 443652
rect 369118 443640 369124 443652
rect 369176 443640 369182 443692
rect 367738 443612 367744 443624
rect 311866 443584 367744 443612
rect 367738 443572 367744 443584
rect 367796 443572 367802 443624
rect 226978 443504 226984 443556
rect 227036 443544 227042 443556
rect 335538 443544 335544 443556
rect 227036 443516 335544 443544
rect 227036 443504 227042 443516
rect 335538 443504 335544 443516
rect 335596 443504 335602 443556
rect 225598 443436 225604 443488
rect 225656 443476 225662 443488
rect 340230 443476 340236 443488
rect 225656 443448 340236 443476
rect 225656 443436 225662 443448
rect 340230 443436 340236 443448
rect 340288 443436 340294 443488
rect 220078 443368 220084 443420
rect 220136 443408 220142 443420
rect 342438 443408 342444 443420
rect 220136 443380 342444 443408
rect 220136 443368 220142 443380
rect 342438 443368 342444 443380
rect 342496 443368 342502 443420
rect 228634 443300 228640 443352
rect 228692 443340 228698 443352
rect 354214 443340 354220 443352
rect 228692 443312 354220 443340
rect 228692 443300 228698 443312
rect 354214 443300 354220 443312
rect 354272 443300 354278 443352
rect 221458 443232 221464 443284
rect 221516 443272 221522 443284
rect 354950 443272 354956 443284
rect 221516 443244 354956 443272
rect 221516 443232 221522 443244
rect 354950 443232 354956 443244
rect 355008 443232 355014 443284
rect 298002 443164 298008 443216
rect 298060 443204 298066 443216
rect 446398 443204 446404 443216
rect 298060 443176 446404 443204
rect 298060 443164 298066 443176
rect 446398 443164 446404 443176
rect 446456 443164 446462 443216
rect 98638 443096 98644 443148
rect 98696 443136 98702 443148
rect 356422 443136 356428 443148
rect 98696 443108 356428 443136
rect 98696 443096 98702 443108
rect 356422 443096 356428 443108
rect 356480 443096 356486 443148
rect 95970 443028 95976 443080
rect 96028 443068 96034 443080
rect 357434 443068 357440 443080
rect 96028 443040 357440 443068
rect 96028 443028 96034 443040
rect 357434 443028 357440 443040
rect 357492 443028 357498 443080
rect 358814 443028 358820 443080
rect 358872 443028 358878 443080
rect 79318 442960 79324 443012
rect 79376 443000 79382 443012
rect 358832 443000 358860 443028
rect 79376 442972 358860 443000
rect 79376 442960 79382 442972
rect 3602 442212 3608 442264
rect 3660 442252 3666 442264
rect 229830 442252 229836 442264
rect 3660 442224 229836 442252
rect 3660 442212 3666 442224
rect 229830 442212 229836 442224
rect 229888 442212 229894 442264
rect 362310 439492 362316 439544
rect 362368 439532 362374 439544
rect 580994 439532 581000 439544
rect 362368 439504 581000 439532
rect 362368 439492 362374 439504
rect 580994 439492 581000 439504
rect 581052 439492 581058 439544
rect 458818 438132 458824 438184
rect 458876 438172 458882 438184
rect 582374 438172 582380 438184
rect 458876 438144 582380 438172
rect 458876 438132 458882 438144
rect 582374 438132 582380 438144
rect 582432 438132 582438 438184
rect 3418 423580 3424 423632
rect 3476 423620 3482 423632
rect 7558 423620 7564 423632
rect 3476 423592 7564 423620
rect 3476 423580 3482 423592
rect 7558 423580 7564 423592
rect 7616 423580 7622 423632
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 226978 411244 226984 411256
rect 3016 411216 226984 411244
rect 3016 411204 3022 411216
rect 226978 411204 226984 411216
rect 227036 411204 227042 411256
rect 3418 410524 3424 410576
rect 3476 410564 3482 410576
rect 229738 410564 229744 410576
rect 3476 410536 229744 410564
rect 3476 410524 3482 410536
rect 229738 410524 229744 410536
rect 229796 410524 229802 410576
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 228634 398800 228640 398812
rect 3384 398772 228640 398800
rect 3384 398760 3390 398772
rect 228634 398760 228640 398772
rect 228692 398760 228698 398812
rect 369118 379448 369124 379500
rect 369176 379488 369182 379500
rect 580166 379488 580172 379500
rect 369176 379460 580172 379488
rect 369176 379448 369182 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3050 372512 3056 372564
rect 3108 372552 3114 372564
rect 228542 372552 228548 372564
rect 3108 372524 228548 372552
rect 3108 372512 3114 372524
rect 228542 372512 228548 372524
rect 228600 372512 228606 372564
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 221458 346372 221464 346384
rect 3384 346344 221464 346372
rect 3384 346332 3390 346344
rect 221458 346332 221464 346344
rect 221516 346332 221522 346384
rect 362218 325592 362224 325644
rect 362276 325632 362282 325644
rect 579890 325632 579896 325644
rect 362276 325604 579896 325632
rect 362276 325592 362282 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 225690 320124 225696 320136
rect 3384 320096 225696 320124
rect 3384 320084 3390 320096
rect 225690 320084 225696 320096
rect 225748 320084 225754 320136
rect 261018 310496 261024 310548
rect 261076 310536 261082 310548
rect 261202 310536 261208 310548
rect 261076 310508 261208 310536
rect 261076 310496 261082 310508
rect 261202 310496 261208 310508
rect 261260 310496 261266 310548
rect 266538 310496 266544 310548
rect 266596 310536 266602 310548
rect 266722 310536 266728 310548
rect 266596 310508 266728 310536
rect 266596 310496 266602 310508
rect 266722 310496 266728 310508
rect 266780 310496 266786 310548
rect 291470 310496 291476 310548
rect 291528 310536 291534 310548
rect 291654 310536 291660 310548
rect 291528 310508 291660 310536
rect 291528 310496 291534 310508
rect 291654 310496 291660 310508
rect 291712 310496 291718 310548
rect 292758 310496 292764 310548
rect 292816 310536 292822 310548
rect 292942 310536 292948 310548
rect 292816 310508 292948 310536
rect 292816 310496 292822 310508
rect 292942 310496 292948 310508
rect 293000 310496 293006 310548
rect 300854 310496 300860 310548
rect 300912 310536 300918 310548
rect 301222 310536 301228 310548
rect 300912 310508 301228 310536
rect 300912 310496 300918 310508
rect 301222 310496 301228 310508
rect 301280 310496 301286 310548
rect 310606 310496 310612 310548
rect 310664 310536 310670 310548
rect 310790 310536 310796 310548
rect 310664 310508 310796 310536
rect 310664 310496 310670 310508
rect 310790 310496 310796 310508
rect 310848 310496 310854 310548
rect 327350 310496 327356 310548
rect 327408 310536 327414 310548
rect 327534 310536 327540 310548
rect 327408 310508 327540 310536
rect 327408 310496 327414 310508
rect 327534 310496 327540 310508
rect 327592 310496 327598 310548
rect 353478 310496 353484 310548
rect 353536 310536 353542 310548
rect 353662 310536 353668 310548
rect 353536 310508 353668 310536
rect 353536 310496 353542 310508
rect 353662 310496 353668 310508
rect 353720 310496 353726 310548
rect 44818 309748 44824 309800
rect 44876 309788 44882 309800
rect 361114 309788 361120 309800
rect 44876 309760 361120 309788
rect 44876 309748 44882 309760
rect 361114 309748 361120 309760
rect 361172 309748 361178 309800
rect 229646 309068 229652 309120
rect 229704 309108 229710 309120
rect 236546 309108 236552 309120
rect 229704 309080 236552 309108
rect 229704 309068 229710 309080
rect 236546 309068 236552 309080
rect 236604 309068 236610 309120
rect 284110 309068 284116 309120
rect 284168 309108 284174 309120
rect 338574 309108 338580 309120
rect 284168 309080 338580 309108
rect 284168 309068 284174 309080
rect 338574 309068 338580 309080
rect 338632 309068 338638 309120
rect 342162 309068 342168 309120
rect 342220 309108 342226 309120
rect 342898 309108 342904 309120
rect 342220 309080 342904 309108
rect 342220 309068 342226 309080
rect 342898 309068 342904 309080
rect 342956 309068 342962 309120
rect 237190 309040 237196 309052
rect 219406 309012 237196 309040
rect 95878 308932 95884 308984
rect 95936 308972 95942 308984
rect 219406 308972 219434 309012
rect 237190 309000 237196 309012
rect 237248 309000 237254 309052
rect 290274 309000 290280 309052
rect 290332 309040 290338 309052
rect 293494 309040 293500 309052
rect 290332 309012 293500 309040
rect 290332 309000 290338 309012
rect 293494 309000 293500 309012
rect 293552 309000 293558 309052
rect 296254 309000 296260 309052
rect 296312 309040 296318 309052
rect 352926 309040 352932 309052
rect 296312 309012 352932 309040
rect 296312 309000 296318 309012
rect 352926 309000 352932 309012
rect 352984 309000 352990 309052
rect 95936 308944 219434 308972
rect 95936 308932 95942 308944
rect 229738 308932 229744 308984
rect 229796 308972 229802 308984
rect 235902 308972 235908 308984
rect 229796 308944 235908 308972
rect 229796 308932 229802 308944
rect 235902 308932 235908 308944
rect 235960 308932 235966 308984
rect 247678 308972 247684 308984
rect 244246 308944 247684 308972
rect 97258 308864 97264 308916
rect 97316 308904 97322 308916
rect 244246 308904 244274 308944
rect 247678 308932 247684 308944
rect 247736 308932 247742 308984
rect 286410 308932 286416 308984
rect 286468 308972 286474 308984
rect 350902 308972 350908 308984
rect 286468 308944 350908 308972
rect 286468 308932 286474 308944
rect 350902 308932 350908 308944
rect 350960 308932 350966 308984
rect 355042 308932 355048 308984
rect 355100 308972 355106 308984
rect 355100 308944 364334 308972
rect 355100 308932 355106 308944
rect 97316 308876 244274 308904
rect 97316 308864 97322 308876
rect 282822 308864 282828 308916
rect 282880 308904 282886 308916
rect 348142 308904 348148 308916
rect 282880 308876 348148 308904
rect 282880 308864 282886 308876
rect 348142 308864 348148 308876
rect 348200 308864 348206 308916
rect 354646 308876 360332 308904
rect 71038 308796 71044 308848
rect 71096 308836 71102 308848
rect 234614 308836 234620 308848
rect 71096 308808 234620 308836
rect 71096 308796 71102 308808
rect 234614 308796 234620 308808
rect 234672 308796 234678 308848
rect 242250 308796 242256 308848
rect 242308 308836 242314 308848
rect 260926 308836 260932 308848
rect 242308 308808 260932 308836
rect 242308 308796 242314 308808
rect 260926 308796 260932 308808
rect 260984 308796 260990 308848
rect 283926 308796 283932 308848
rect 283984 308836 283990 308848
rect 352006 308836 352012 308848
rect 283984 308808 352012 308836
rect 283984 308796 283990 308808
rect 352006 308796 352012 308808
rect 352064 308796 352070 308848
rect 64138 308728 64144 308780
rect 64196 308768 64202 308780
rect 232866 308768 232872 308780
rect 64196 308740 232872 308768
rect 64196 308728 64202 308740
rect 232866 308728 232872 308740
rect 232924 308728 232930 308780
rect 235810 308728 235816 308780
rect 235868 308768 235874 308780
rect 243722 308768 243728 308780
rect 235868 308740 243728 308768
rect 235868 308728 235874 308740
rect 243722 308728 243728 308740
rect 243780 308728 243786 308780
rect 275554 308728 275560 308780
rect 275612 308768 275618 308780
rect 279878 308768 279884 308780
rect 275612 308740 279884 308768
rect 275612 308728 275618 308740
rect 279878 308728 279884 308740
rect 279936 308728 279942 308780
rect 285582 308728 285588 308780
rect 285640 308768 285646 308780
rect 354030 308768 354036 308780
rect 285640 308740 354036 308768
rect 285640 308728 285646 308740
rect 354030 308728 354036 308740
rect 354088 308728 354094 308780
rect 46198 308660 46204 308712
rect 46256 308700 46262 308712
rect 229646 308700 229652 308712
rect 46256 308672 229652 308700
rect 46256 308660 46262 308672
rect 229646 308660 229652 308672
rect 229704 308660 229710 308712
rect 257338 308660 257344 308712
rect 257396 308700 257402 308712
rect 277026 308700 277032 308712
rect 257396 308672 277032 308700
rect 257396 308660 257402 308672
rect 277026 308660 277032 308672
rect 277084 308660 277090 308712
rect 287698 308660 287704 308712
rect 287756 308700 287762 308712
rect 348786 308700 348792 308712
rect 287756 308672 348792 308700
rect 287756 308660 287762 308672
rect 348786 308660 348792 308672
rect 348844 308660 348850 308712
rect 354398 308660 354404 308712
rect 354456 308700 354462 308712
rect 354646 308700 354674 308876
rect 355686 308728 355692 308780
rect 355744 308768 355750 308780
rect 355744 308740 360240 308768
rect 355744 308728 355750 308740
rect 354456 308672 354674 308700
rect 354456 308660 354462 308672
rect 31754 308592 31760 308644
rect 31812 308632 31818 308644
rect 229738 308632 229744 308644
rect 31812 308604 229744 308632
rect 31812 308592 31818 308604
rect 229738 308592 229744 308604
rect 229796 308592 229802 308644
rect 243722 308592 243728 308644
rect 243780 308632 243786 308644
rect 251174 308632 251180 308644
rect 243780 308604 251180 308632
rect 243780 308592 243786 308604
rect 251174 308592 251180 308604
rect 251232 308592 251238 308644
rect 253566 308592 253572 308644
rect 253624 308632 253630 308644
rect 254394 308632 254400 308644
rect 253624 308604 254400 308632
rect 253624 308592 253630 308604
rect 254394 308592 254400 308604
rect 254452 308592 254458 308644
rect 279878 308592 279884 308644
rect 279936 308632 279942 308644
rect 349430 308632 349436 308644
rect 279936 308604 349436 308632
rect 279936 308592 279942 308604
rect 349430 308592 349436 308604
rect 349488 308592 349494 308644
rect 356238 308592 356244 308644
rect 356296 308632 356302 308644
rect 356422 308632 356428 308644
rect 356296 308604 356428 308632
rect 356296 308592 356302 308604
rect 356422 308592 356428 308604
rect 356480 308592 356486 308644
rect 358998 308592 359004 308644
rect 359056 308632 359062 308644
rect 359274 308632 359280 308644
rect 359056 308604 359280 308632
rect 359056 308592 359062 308604
rect 359274 308592 359280 308604
rect 359332 308592 359338 308644
rect 360212 308632 360240 308740
rect 360304 308700 360332 308876
rect 364306 308768 364334 308944
rect 438026 308768 438032 308780
rect 364306 308740 438032 308768
rect 438026 308728 438032 308740
rect 438084 308728 438090 308780
rect 436830 308700 436836 308712
rect 360304 308672 436836 308700
rect 436830 308660 436836 308672
rect 436888 308660 436894 308712
rect 439498 308632 439504 308644
rect 360212 308604 439504 308632
rect 439498 308592 439504 308604
rect 439556 308592 439562 308644
rect 39298 308524 39304 308576
rect 39356 308564 39362 308576
rect 232038 308564 232044 308576
rect 39356 308536 232044 308564
rect 39356 308524 39362 308536
rect 232038 308524 232044 308536
rect 232096 308524 232102 308576
rect 249058 308524 249064 308576
rect 249116 308564 249122 308576
rect 347682 308564 347688 308576
rect 249116 308536 347688 308564
rect 249116 308524 249122 308536
rect 347682 308524 347688 308536
rect 347740 308524 347746 308576
rect 353754 308524 353760 308576
rect 353812 308564 353818 308576
rect 439590 308564 439596 308576
rect 353812 308536 439596 308564
rect 353812 308524 353818 308536
rect 439590 308524 439596 308536
rect 439648 308524 439654 308576
rect 27614 308456 27620 308508
rect 27672 308496 27678 308508
rect 235258 308496 235264 308508
rect 27672 308468 235264 308496
rect 27672 308456 27678 308468
rect 235258 308456 235264 308468
rect 235316 308456 235322 308508
rect 236822 308456 236828 308508
rect 236880 308496 236886 308508
rect 246390 308496 246396 308508
rect 236880 308468 246396 308496
rect 236880 308456 236886 308468
rect 246390 308456 246396 308468
rect 246448 308456 246454 308508
rect 247678 308456 247684 308508
rect 247736 308496 247742 308508
rect 348970 308496 348976 308508
rect 247736 308468 348976 308496
rect 247736 308456 247742 308468
rect 348970 308456 348976 308468
rect 349028 308456 349034 308508
rect 353110 308456 353116 308508
rect 353168 308496 353174 308508
rect 438118 308496 438124 308508
rect 353168 308468 438124 308496
rect 353168 308456 353174 308468
rect 438118 308456 438124 308468
rect 438176 308456 438182 308508
rect 23474 308388 23480 308440
rect 23532 308428 23538 308440
rect 234430 308428 234436 308440
rect 23532 308400 234436 308428
rect 23532 308388 23538 308400
rect 234430 308388 234436 308400
rect 234488 308388 234494 308440
rect 238018 308388 238024 308440
rect 238076 308428 238082 308440
rect 238076 308400 331214 308428
rect 238076 308388 238082 308400
rect 282638 308320 282644 308372
rect 282696 308360 282702 308372
rect 283650 308360 283656 308372
rect 282696 308332 283656 308360
rect 282696 308320 282702 308332
rect 283650 308320 283656 308332
rect 283708 308320 283714 308372
rect 331186 308360 331214 308400
rect 340874 308388 340880 308440
rect 340932 308428 340938 308440
rect 341886 308428 341892 308440
rect 340932 308400 341892 308428
rect 340932 308388 340938 308400
rect 341886 308388 341892 308400
rect 341944 308388 341950 308440
rect 342530 308388 342536 308440
rect 342588 308428 342594 308440
rect 343174 308428 343180 308440
rect 342588 308400 343180 308428
rect 342588 308388 342594 308400
rect 343174 308388 343180 308400
rect 343232 308388 343238 308440
rect 343634 308388 343640 308440
rect 343692 308428 343698 308440
rect 343910 308428 343916 308440
rect 343692 308400 343916 308428
rect 343692 308388 343698 308400
rect 343910 308388 343916 308400
rect 343968 308388 343974 308440
rect 345198 308388 345204 308440
rect 345256 308428 345262 308440
rect 345934 308428 345940 308440
rect 345256 308400 345940 308428
rect 345256 308388 345262 308400
rect 345934 308388 345940 308400
rect 345992 308388 345998 308440
rect 346578 308388 346584 308440
rect 346636 308428 346642 308440
rect 346854 308428 346860 308440
rect 346636 308400 346860 308428
rect 346636 308388 346642 308400
rect 346854 308388 346860 308400
rect 346912 308388 346918 308440
rect 349338 308388 349344 308440
rect 349396 308428 349402 308440
rect 350074 308428 350080 308440
rect 349396 308400 350080 308428
rect 349396 308388 349402 308400
rect 350074 308388 350080 308400
rect 350132 308388 350138 308440
rect 352466 308388 352472 308440
rect 352524 308428 352530 308440
rect 440510 308428 440516 308440
rect 352524 308400 440516 308428
rect 352524 308388 352530 308400
rect 440510 308388 440516 308400
rect 440568 308388 440574 308440
rect 331186 308332 345014 308360
rect 337470 308292 337476 308304
rect 283852 308264 337476 308292
rect 250438 308184 250444 308236
rect 250496 308224 250502 308236
rect 252646 308224 252652 308236
rect 250496 308196 252652 308224
rect 250496 308184 250502 308196
rect 252646 308184 252652 308196
rect 252704 308184 252710 308236
rect 281442 308184 281448 308236
rect 281500 308224 281506 308236
rect 283742 308224 283748 308236
rect 281500 308196 283748 308224
rect 281500 308184 281506 308196
rect 283742 308184 283748 308196
rect 283800 308184 283806 308236
rect 247586 308116 247592 308168
rect 247644 308156 247650 308168
rect 252278 308156 252284 308168
rect 247644 308128 252284 308156
rect 247644 308116 247650 308128
rect 252278 308116 252284 308128
rect 252336 308116 252342 308168
rect 243630 308048 243636 308100
rect 243688 308088 243694 308100
rect 250070 308088 250076 308100
rect 243688 308060 250076 308088
rect 243688 308048 243694 308060
rect 250070 308048 250076 308060
rect 250128 308048 250134 308100
rect 252646 308048 252652 308100
rect 252704 308088 252710 308100
rect 253290 308088 253296 308100
rect 252704 308060 253296 308088
rect 252704 308048 252710 308060
rect 253290 308048 253296 308060
rect 253348 308048 253354 308100
rect 283742 308048 283748 308100
rect 283800 308088 283806 308100
rect 283852 308088 283880 308264
rect 337470 308252 337476 308264
rect 337528 308252 337534 308304
rect 341150 308252 341156 308304
rect 341208 308292 341214 308304
rect 341794 308292 341800 308304
rect 341208 308264 341800 308292
rect 341208 308252 341214 308264
rect 341794 308252 341800 308264
rect 341852 308252 341858 308304
rect 342622 308252 342628 308304
rect 342680 308292 342686 308304
rect 343542 308292 343548 308304
rect 342680 308264 343548 308292
rect 342680 308252 342686 308264
rect 343542 308252 343548 308264
rect 343600 308252 343606 308304
rect 320174 308184 320180 308236
rect 320232 308224 320238 308236
rect 320726 308224 320732 308236
rect 320232 308196 320732 308224
rect 320232 308184 320238 308196
rect 320726 308184 320732 308196
rect 320784 308184 320790 308236
rect 342346 308184 342352 308236
rect 342404 308224 342410 308236
rect 343082 308224 343088 308236
rect 342404 308196 343088 308224
rect 342404 308184 342410 308196
rect 343082 308184 343088 308196
rect 343140 308184 343146 308236
rect 344986 308224 345014 308332
rect 345106 308320 345112 308372
rect 345164 308360 345170 308372
rect 345566 308360 345572 308372
rect 345164 308332 345572 308360
rect 345164 308320 345170 308332
rect 345566 308320 345572 308332
rect 345624 308320 345630 308372
rect 346670 308320 346676 308372
rect 346728 308360 346734 308372
rect 347222 308360 347228 308372
rect 346728 308332 347228 308360
rect 346728 308320 346734 308332
rect 347222 308320 347228 308332
rect 347280 308320 347286 308372
rect 354674 308320 354680 308372
rect 354732 308360 354738 308372
rect 354858 308360 354864 308372
rect 354732 308332 354864 308360
rect 354732 308320 354738 308332
rect 354858 308320 354864 308332
rect 354916 308320 354922 308372
rect 356146 308320 356152 308372
rect 356204 308360 356210 308372
rect 356790 308360 356796 308372
rect 356204 308332 356796 308360
rect 356204 308320 356210 308332
rect 356790 308320 356796 308332
rect 356848 308320 356854 308372
rect 357526 308320 357532 308372
rect 357584 308360 357590 308372
rect 358078 308360 358084 308372
rect 357584 308332 358084 308360
rect 357584 308320 357590 308332
rect 358078 308320 358084 308332
rect 358136 308320 358142 308372
rect 345290 308252 345296 308304
rect 345348 308292 345354 308304
rect 345474 308292 345480 308304
rect 345348 308264 345480 308292
rect 345348 308252 345354 308264
rect 345474 308252 345480 308264
rect 345532 308252 345538 308304
rect 356054 308252 356060 308304
rect 356112 308292 356118 308304
rect 357250 308292 357256 308304
rect 356112 308264 357256 308292
rect 356112 308252 356118 308264
rect 357250 308252 357256 308264
rect 357308 308252 357314 308304
rect 357710 308252 357716 308304
rect 357768 308292 357774 308304
rect 358170 308292 358176 308304
rect 357768 308264 358176 308292
rect 357768 308252 357774 308264
rect 358170 308252 358176 308264
rect 358228 308252 358234 308304
rect 359182 308252 359188 308304
rect 359240 308292 359246 308304
rect 359826 308292 359832 308304
rect 359240 308264 359832 308292
rect 359240 308252 359246 308264
rect 359826 308252 359832 308264
rect 359884 308252 359890 308304
rect 360194 308252 360200 308304
rect 360252 308292 360258 308304
rect 360470 308292 360476 308304
rect 360252 308264 360476 308292
rect 360252 308252 360258 308264
rect 360470 308252 360476 308264
rect 360528 308252 360534 308304
rect 350258 308224 350264 308236
rect 344986 308196 350264 308224
rect 350258 308184 350264 308196
rect 350316 308184 350322 308236
rect 357618 308184 357624 308236
rect 357676 308224 357682 308236
rect 358538 308224 358544 308236
rect 357676 308196 358544 308224
rect 357676 308184 357682 308196
rect 358538 308184 358544 308196
rect 358596 308184 358602 308236
rect 359090 308184 359096 308236
rect 359148 308224 359154 308236
rect 359918 308224 359924 308236
rect 359148 308196 359924 308224
rect 359148 308184 359154 308196
rect 359918 308184 359924 308196
rect 359976 308184 359982 308236
rect 337654 308156 337660 308168
rect 302206 308128 337660 308156
rect 283800 308060 283880 308088
rect 283800 308048 283806 308060
rect 284386 308048 284392 308100
rect 284444 308088 284450 308100
rect 293218 308088 293224 308100
rect 284444 308060 293224 308088
rect 284444 308048 284450 308060
rect 293218 308048 293224 308060
rect 293276 308048 293282 308100
rect 246390 307980 246396 308032
rect 246448 308020 246454 308032
rect 250254 308020 250260 308032
rect 246448 307992 250260 308020
rect 246448 307980 246454 307992
rect 250254 307980 250260 307992
rect 250312 307980 250318 308032
rect 283558 307980 283564 308032
rect 283616 308020 283622 308032
rect 285214 308020 285220 308032
rect 283616 307992 285220 308020
rect 283616 307980 283622 307992
rect 285214 307980 285220 307992
rect 285272 307980 285278 308032
rect 246850 307912 246856 307964
rect 246908 307952 246914 307964
rect 249886 307952 249892 307964
rect 246908 307924 249892 307952
rect 246908 307912 246914 307924
rect 249886 307912 249892 307924
rect 249944 307912 249950 307964
rect 261202 307912 261208 307964
rect 261260 307952 261266 307964
rect 261662 307952 261668 307964
rect 261260 307924 261668 307952
rect 261260 307912 261266 307924
rect 261662 307912 261668 307924
rect 261720 307912 261726 307964
rect 274082 307912 274088 307964
rect 274140 307952 274146 307964
rect 279418 307952 279424 307964
rect 274140 307924 279424 307952
rect 274140 307912 274146 307924
rect 279418 307912 279424 307924
rect 279476 307912 279482 307964
rect 279786 307912 279792 307964
rect 279844 307952 279850 307964
rect 287698 307952 287704 307964
rect 279844 307924 287704 307952
rect 279844 307912 279850 307924
rect 287698 307912 287704 307924
rect 287756 307912 287762 307964
rect 291010 307912 291016 307964
rect 291068 307952 291074 307964
rect 302206 307952 302234 308128
rect 337654 308116 337660 308128
rect 337712 308116 337718 308168
rect 345290 308116 345296 308168
rect 345348 308156 345354 308168
rect 346118 308156 346124 308168
rect 345348 308128 346124 308156
rect 345348 308116 345354 308128
rect 346118 308116 346124 308128
rect 346176 308116 346182 308168
rect 350810 308116 350816 308168
rect 350868 308156 350874 308168
rect 351454 308156 351460 308168
rect 350868 308128 351460 308156
rect 350868 308116 350874 308128
rect 351454 308116 351460 308128
rect 351512 308116 351518 308168
rect 354766 308116 354772 308168
rect 354824 308156 354830 308168
rect 355502 308156 355508 308168
rect 354824 308128 355508 308156
rect 354824 308116 354830 308128
rect 355502 308116 355508 308128
rect 355560 308116 355566 308168
rect 358814 308116 358820 308168
rect 358872 308156 358878 308168
rect 359458 308156 359464 308168
rect 358872 308128 359464 308156
rect 358872 308116 358878 308128
rect 359458 308116 359464 308128
rect 359516 308116 359522 308168
rect 350626 308048 350632 308100
rect 350684 308088 350690 308100
rect 351362 308088 351368 308100
rect 350684 308060 351368 308088
rect 350684 308048 350690 308060
rect 351362 308048 351368 308060
rect 351420 308048 351426 308100
rect 359274 308048 359280 308100
rect 359332 308048 359338 308100
rect 291068 307924 302234 307952
rect 291068 307912 291074 307924
rect 240870 307844 240876 307896
rect 240928 307884 240934 307896
rect 240928 307856 244274 307884
rect 240928 307844 240934 307856
rect 229738 307776 229744 307828
rect 229796 307816 229802 307828
rect 230934 307816 230940 307828
rect 229796 307788 230940 307816
rect 229796 307776 229802 307788
rect 230934 307776 230940 307788
rect 230992 307776 230998 307828
rect 236730 307776 236736 307828
rect 236788 307816 236794 307828
rect 238110 307816 238116 307828
rect 236788 307788 238116 307816
rect 236788 307776 236794 307788
rect 238110 307776 238116 307788
rect 238168 307776 238174 307828
rect 239766 307776 239772 307828
rect 239824 307816 239830 307828
rect 241146 307816 241152 307828
rect 239824 307788 241152 307816
rect 239824 307776 239830 307788
rect 241146 307776 241152 307788
rect 241204 307776 241210 307828
rect 242158 307776 242164 307828
rect 242216 307816 242222 307828
rect 242894 307816 242900 307828
rect 242216 307788 242900 307816
rect 242216 307776 242222 307788
rect 242894 307776 242900 307788
rect 242952 307776 242958 307828
rect 244246 307816 244274 307856
rect 246298 307844 246304 307896
rect 246356 307884 246362 307896
rect 248966 307884 248972 307896
rect 246356 307856 248972 307884
rect 246356 307844 246362 307856
rect 248966 307844 248972 307856
rect 249024 307844 249030 307896
rect 253382 307844 253388 307896
rect 253440 307884 253446 307896
rect 259638 307884 259644 307896
rect 253440 307856 259644 307884
rect 253440 307844 253446 307856
rect 259638 307844 259644 307856
rect 259696 307844 259702 307896
rect 260098 307844 260104 307896
rect 260156 307884 260162 307896
rect 262858 307884 262864 307896
rect 260156 307856 262864 307884
rect 260156 307844 260162 307856
rect 262858 307844 262864 307856
rect 262916 307844 262922 307896
rect 268470 307844 268476 307896
rect 268528 307884 268534 307896
rect 275738 307884 275744 307896
rect 268528 307856 275744 307884
rect 268528 307844 268534 307856
rect 275738 307844 275744 307856
rect 275796 307844 275802 307896
rect 278866 307844 278872 307896
rect 278924 307884 278930 307896
rect 281350 307884 281356 307896
rect 278924 307856 281356 307884
rect 278924 307844 278930 307856
rect 281350 307844 281356 307856
rect 281408 307844 281414 307896
rect 284662 307844 284668 307896
rect 284720 307884 284726 307896
rect 286318 307884 286324 307896
rect 284720 307856 286324 307884
rect 284720 307844 284726 307856
rect 286318 307844 286324 307856
rect 286376 307844 286382 307896
rect 293954 307844 293960 307896
rect 294012 307884 294018 307896
rect 295794 307884 295800 307896
rect 294012 307856 295800 307884
rect 294012 307844 294018 307856
rect 295794 307844 295800 307856
rect 295852 307844 295858 307896
rect 317506 307844 317512 307896
rect 317564 307884 317570 307896
rect 320818 307884 320824 307896
rect 317564 307856 320824 307884
rect 317564 307844 317570 307856
rect 320818 307844 320824 307856
rect 320876 307844 320882 307896
rect 334250 307844 334256 307896
rect 334308 307884 334314 307896
rect 334802 307884 334808 307896
rect 334308 307856 334808 307884
rect 334308 307844 334314 307856
rect 334802 307844 334808 307856
rect 334860 307844 334866 307896
rect 359292 307884 359320 308048
rect 359366 307884 359372 307896
rect 359292 307856 359372 307884
rect 359366 307844 359372 307856
rect 359424 307844 359430 307896
rect 247678 307816 247684 307828
rect 244246 307788 247684 307816
rect 247678 307776 247684 307788
rect 247736 307776 247742 307828
rect 247770 307776 247776 307828
rect 247828 307816 247834 307828
rect 248506 307816 248512 307828
rect 247828 307788 248512 307816
rect 247828 307776 247834 307788
rect 248506 307776 248512 307788
rect 248564 307776 248570 307828
rect 253290 307776 253296 307828
rect 253348 307816 253354 307828
rect 253566 307816 253572 307828
rect 253348 307788 253572 307816
rect 253348 307776 253354 307788
rect 253566 307776 253572 307788
rect 253624 307776 253630 307828
rect 254946 307776 254952 307828
rect 255004 307816 255010 307828
rect 255682 307816 255688 307828
rect 255004 307788 255688 307816
rect 255004 307776 255010 307788
rect 255682 307776 255688 307788
rect 255740 307776 255746 307828
rect 256234 307776 256240 307828
rect 256292 307816 256298 307828
rect 258350 307816 258356 307828
rect 256292 307788 258356 307816
rect 256292 307776 256298 307788
rect 258350 307776 258356 307788
rect 258408 307776 258414 307828
rect 261662 307776 261668 307828
rect 261720 307816 261726 307828
rect 262214 307816 262220 307828
rect 261720 307788 262220 307816
rect 261720 307776 261726 307788
rect 262214 307776 262220 307788
rect 262272 307776 262278 307828
rect 265618 307776 265624 307828
rect 265676 307816 265682 307828
rect 266814 307816 266820 307828
rect 265676 307788 266820 307816
rect 265676 307776 265682 307788
rect 266814 307776 266820 307788
rect 266872 307776 266878 307828
rect 269758 307776 269764 307828
rect 269816 307816 269822 307828
rect 272058 307816 272064 307828
rect 269816 307788 272064 307816
rect 269816 307776 269822 307788
rect 272058 307776 272064 307788
rect 272116 307776 272122 307828
rect 278038 307776 278044 307828
rect 278096 307816 278102 307828
rect 278958 307816 278964 307828
rect 278096 307788 278964 307816
rect 278096 307776 278102 307788
rect 278958 307776 278964 307788
rect 279016 307776 279022 307828
rect 279694 307776 279700 307828
rect 279752 307816 279758 307828
rect 281166 307816 281172 307828
rect 279752 307788 281172 307816
rect 279752 307776 279758 307788
rect 281166 307776 281172 307788
rect 281224 307776 281230 307828
rect 284018 307776 284024 307828
rect 284076 307816 284082 307828
rect 284938 307816 284944 307828
rect 284076 307788 284944 307816
rect 284076 307776 284082 307788
rect 284938 307776 284944 307788
rect 284996 307776 285002 307828
rect 286778 307776 286784 307828
rect 286836 307816 286842 307828
rect 289078 307816 289084 307828
rect 286836 307788 289084 307816
rect 286836 307776 286842 307788
rect 289078 307776 289084 307788
rect 289136 307776 289142 307828
rect 292666 307776 292672 307828
rect 292724 307816 292730 307828
rect 294506 307816 294512 307828
rect 292724 307788 294512 307816
rect 292724 307776 292730 307788
rect 294506 307776 294512 307788
rect 294564 307776 294570 307828
rect 295242 307776 295248 307828
rect 295300 307816 295306 307828
rect 296070 307816 296076 307828
rect 295300 307788 296076 307816
rect 295300 307776 295306 307788
rect 296070 307776 296076 307788
rect 296128 307776 296134 307828
rect 314838 307776 314844 307828
rect 314896 307816 314902 307828
rect 318058 307816 318064 307828
rect 314896 307788 318064 307816
rect 314896 307776 314902 307788
rect 318058 307776 318064 307788
rect 318116 307776 318122 307828
rect 343634 307232 343640 307284
rect 343692 307272 343698 307284
rect 344646 307272 344652 307284
rect 343692 307244 344652 307272
rect 343692 307232 343698 307244
rect 344646 307232 344652 307244
rect 344704 307232 344710 307284
rect 68278 307164 68284 307216
rect 68336 307204 68342 307216
rect 241790 307204 241796 307216
rect 68336 307176 241796 307204
rect 68336 307164 68342 307176
rect 241790 307164 241796 307176
rect 241848 307164 241854 307216
rect 334618 307164 334624 307216
rect 334676 307204 334682 307216
rect 445018 307204 445024 307216
rect 334676 307176 445024 307204
rect 334676 307164 334682 307176
rect 445018 307164 445024 307176
rect 445076 307164 445082 307216
rect 57974 307096 57980 307148
rect 58032 307136 58038 307148
rect 240686 307136 240692 307148
rect 58032 307108 240692 307136
rect 58032 307096 58038 307108
rect 240686 307096 240692 307108
rect 240744 307096 240750 307148
rect 318334 307096 318340 307148
rect 318392 307136 318398 307148
rect 462958 307136 462964 307148
rect 318392 307108 462964 307136
rect 318392 307096 318398 307108
rect 462958 307096 462964 307108
rect 463016 307096 463022 307148
rect 25498 307028 25504 307080
rect 25556 307068 25562 307080
rect 230106 307068 230112 307080
rect 25556 307040 230112 307068
rect 25556 307028 25562 307040
rect 230106 307028 230112 307040
rect 230164 307028 230170 307080
rect 238018 307028 238024 307080
rect 238076 307068 238082 307080
rect 252922 307068 252928 307080
rect 238076 307040 252928 307068
rect 238076 307028 238082 307040
rect 252922 307028 252928 307040
rect 252980 307028 252986 307080
rect 264238 307028 264244 307080
rect 264296 307068 264302 307080
rect 274634 307068 274640 307080
rect 264296 307040 274640 307068
rect 264296 307028 264302 307040
rect 274634 307028 274640 307040
rect 274692 307028 274698 307080
rect 322198 307028 322204 307080
rect 322256 307068 322262 307080
rect 500218 307068 500224 307080
rect 322256 307040 500224 307068
rect 322256 307028 322262 307040
rect 500218 307028 500224 307040
rect 500276 307028 500282 307080
rect 257062 306960 257068 307012
rect 257120 306960 257126 307012
rect 268102 306960 268108 307012
rect 268160 306960 268166 307012
rect 287238 306960 287244 307012
rect 287296 306960 287302 307012
rect 257080 306796 257108 306960
rect 257154 306796 257160 306808
rect 257080 306768 257160 306796
rect 257154 306756 257160 306768
rect 257212 306756 257218 306808
rect 268120 306796 268148 306960
rect 268194 306796 268200 306808
rect 268120 306768 268200 306796
rect 268194 306756 268200 306768
rect 268252 306756 268258 306808
rect 287256 306796 287284 306960
rect 287330 306796 287336 306808
rect 287256 306768 287336 306796
rect 287330 306756 287336 306768
rect 287388 306756 287394 306808
rect 233510 306688 233516 306740
rect 233568 306688 233574 306740
rect 259822 306688 259828 306740
rect 259880 306688 259886 306740
rect 233528 306536 233556 306688
rect 233510 306484 233516 306536
rect 233568 306484 233574 306536
rect 238754 306484 238760 306536
rect 238812 306524 238818 306536
rect 239122 306524 239128 306536
rect 238812 306496 239128 306524
rect 238812 306484 238818 306496
rect 239122 306484 239128 306496
rect 239180 306484 239186 306536
rect 245654 306484 245660 306536
rect 245712 306524 245718 306536
rect 245930 306524 245936 306536
rect 245712 306496 245936 306524
rect 245712 306484 245718 306496
rect 245930 306484 245936 306496
rect 245988 306484 245994 306536
rect 259840 306468 259868 306688
rect 320266 306620 320272 306672
rect 320324 306660 320330 306672
rect 321094 306660 321100 306672
rect 320324 306632 321100 306660
rect 320324 306620 320330 306632
rect 321094 306620 321100 306632
rect 321152 306620 321158 306672
rect 303798 306552 303804 306604
rect 303856 306592 303862 306604
rect 304350 306592 304356 306604
rect 303856 306564 304356 306592
rect 303856 306552 303862 306564
rect 304350 306552 304356 306564
rect 304408 306552 304414 306604
rect 325786 306552 325792 306604
rect 325844 306592 325850 306604
rect 326798 306592 326804 306604
rect 325844 306564 326804 306592
rect 325844 306552 325850 306564
rect 326798 306552 326804 306564
rect 326856 306552 326862 306604
rect 350718 306552 350724 306604
rect 350776 306592 350782 306604
rect 351822 306592 351828 306604
rect 350776 306564 351828 306592
rect 350776 306552 350782 306564
rect 351822 306552 351828 306564
rect 351880 306552 351886 306604
rect 287146 306484 287152 306536
rect 287204 306524 287210 306536
rect 287422 306524 287428 306536
rect 287204 306496 287428 306524
rect 287204 306484 287210 306496
rect 287422 306484 287428 306496
rect 287480 306484 287486 306536
rect 292666 306484 292672 306536
rect 292724 306524 292730 306536
rect 293770 306524 293776 306536
rect 292724 306496 293776 306524
rect 292724 306484 292730 306496
rect 293770 306484 293776 306496
rect 293828 306484 293834 306536
rect 294046 306484 294052 306536
rect 294104 306524 294110 306536
rect 295058 306524 295064 306536
rect 294104 306496 295064 306524
rect 294104 306484 294110 306496
rect 295058 306484 295064 306496
rect 295116 306484 295122 306536
rect 295426 306484 295432 306536
rect 295484 306524 295490 306536
rect 296162 306524 296168 306536
rect 295484 306496 296168 306524
rect 295484 306484 295490 306496
rect 296162 306484 296168 306496
rect 296220 306484 296226 306536
rect 299566 306484 299572 306536
rect 299624 306524 299630 306536
rect 300118 306524 300124 306536
rect 299624 306496 300124 306524
rect 299624 306484 299630 306496
rect 300118 306484 300124 306496
rect 300176 306484 300182 306536
rect 302418 306484 302424 306536
rect 302476 306524 302482 306536
rect 303338 306524 303344 306536
rect 302476 306496 303344 306524
rect 302476 306484 302482 306496
rect 303338 306484 303344 306496
rect 303396 306484 303402 306536
rect 313734 306484 313740 306536
rect 313792 306524 313798 306536
rect 313918 306524 313924 306536
rect 313792 306496 313924 306524
rect 313792 306484 313798 306496
rect 313918 306484 313924 306496
rect 313976 306484 313982 306536
rect 316126 306484 316132 306536
rect 316184 306524 316190 306536
rect 317230 306524 317236 306536
rect 316184 306496 317236 306524
rect 316184 306484 316190 306496
rect 317230 306484 317236 306496
rect 317288 306484 317294 306536
rect 320266 306484 320272 306536
rect 320324 306524 320330 306536
rect 321002 306524 321008 306536
rect 320324 306496 321008 306524
rect 320324 306484 320330 306496
rect 321002 306484 321008 306496
rect 321060 306484 321066 306536
rect 325878 306484 325884 306536
rect 325936 306524 325942 306536
rect 326246 306524 326252 306536
rect 325936 306496 326252 306524
rect 325936 306484 325942 306496
rect 326246 306484 326252 306496
rect 326304 306484 326310 306536
rect 327166 306484 327172 306536
rect 327224 306524 327230 306536
rect 328178 306524 328184 306536
rect 327224 306496 328184 306524
rect 327224 306484 327230 306496
rect 328178 306484 328184 306496
rect 328236 306484 328242 306536
rect 331214 306484 331220 306536
rect 331272 306524 331278 306536
rect 331766 306524 331772 306536
rect 331272 306496 331772 306524
rect 331272 306484 331278 306496
rect 331766 306484 331772 306496
rect 331824 306484 331830 306536
rect 333974 306484 333980 306536
rect 334032 306524 334038 306536
rect 334526 306524 334532 306536
rect 334032 306496 334532 306524
rect 334032 306484 334038 306496
rect 334526 306484 334532 306496
rect 334584 306484 334590 306536
rect 234706 306416 234712 306468
rect 234764 306456 234770 306468
rect 235350 306456 235356 306468
rect 234764 306428 235356 306456
rect 234764 306416 234770 306428
rect 235350 306416 235356 306428
rect 235408 306416 235414 306468
rect 239398 306456 239404 306468
rect 238864 306428 239404 306456
rect 232038 306348 232044 306400
rect 232096 306388 232102 306400
rect 232958 306388 232964 306400
rect 232096 306360 232964 306388
rect 232096 306348 232102 306360
rect 232958 306348 232964 306360
rect 233016 306348 233022 306400
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 225598 306320 225604 306332
rect 3384 306292 225604 306320
rect 3384 306280 3390 306292
rect 225598 306280 225604 306292
rect 225656 306280 225662 306332
rect 229186 306280 229192 306332
rect 229244 306320 229250 306332
rect 230290 306320 230296 306332
rect 229244 306292 230296 306320
rect 229244 306280 229250 306292
rect 230290 306280 230296 306292
rect 230348 306280 230354 306332
rect 231946 306280 231952 306332
rect 232004 306320 232010 306332
rect 232498 306320 232504 306332
rect 232004 306292 232504 306320
rect 232004 306280 232010 306292
rect 232498 306280 232504 306292
rect 232556 306280 232562 306332
rect 236178 306280 236184 306332
rect 236236 306320 236242 306332
rect 237006 306320 237012 306332
rect 236236 306292 237012 306320
rect 236236 306280 236242 306292
rect 237006 306280 237012 306292
rect 237064 306280 237070 306332
rect 238864 306264 238892 306428
rect 239398 306416 239404 306428
rect 239456 306416 239462 306468
rect 245838 306416 245844 306468
rect 245896 306456 245902 306468
rect 246574 306456 246580 306468
rect 245896 306428 246580 306456
rect 245896 306416 245902 306428
rect 246574 306416 246580 306428
rect 246632 306416 246638 306468
rect 259822 306416 259828 306468
rect 259880 306416 259886 306468
rect 272058 306416 272064 306468
rect 272116 306456 272122 306468
rect 272886 306456 272892 306468
rect 272116 306428 272892 306456
rect 272116 306416 272122 306428
rect 272886 306416 272892 306428
rect 272944 306416 272950 306468
rect 273438 306416 273444 306468
rect 273496 306456 273502 306468
rect 273622 306456 273628 306468
rect 273496 306428 273628 306456
rect 273496 306416 273502 306428
rect 273622 306416 273628 306428
rect 273680 306416 273686 306468
rect 281626 306416 281632 306468
rect 281684 306456 281690 306468
rect 282178 306456 282184 306468
rect 281684 306428 282184 306456
rect 281684 306416 281690 306428
rect 282178 306416 282184 306428
rect 282236 306416 282242 306468
rect 285674 306416 285680 306468
rect 285732 306456 285738 306468
rect 286594 306456 286600 306468
rect 285732 306428 286600 306456
rect 285732 306416 285738 306428
rect 286594 306416 286600 306428
rect 286652 306416 286658 306468
rect 287054 306416 287060 306468
rect 287112 306456 287118 306468
rect 287606 306456 287612 306468
rect 287112 306428 287612 306456
rect 287112 306416 287118 306428
rect 287606 306416 287612 306428
rect 287664 306416 287670 306468
rect 288526 306416 288532 306468
rect 288584 306456 288590 306468
rect 288802 306456 288808 306468
rect 288584 306428 288808 306456
rect 288584 306416 288590 306428
rect 288802 306416 288808 306428
rect 288860 306416 288866 306468
rect 292574 306416 292580 306468
rect 292632 306456 292638 306468
rect 293310 306456 293316 306468
rect 292632 306428 293316 306456
rect 292632 306416 292638 306428
rect 293310 306416 293316 306428
rect 293368 306416 293374 306468
rect 293954 306416 293960 306468
rect 294012 306456 294018 306468
rect 294414 306456 294420 306468
rect 294012 306428 294420 306456
rect 294012 306416 294018 306428
rect 294414 306416 294420 306428
rect 294472 306416 294478 306468
rect 295610 306416 295616 306468
rect 295668 306456 295674 306468
rect 296346 306456 296352 306468
rect 295668 306428 296352 306456
rect 295668 306416 295674 306428
rect 296346 306416 296352 306428
rect 296404 306416 296410 306468
rect 299474 306416 299480 306468
rect 299532 306456 299538 306468
rect 300026 306456 300032 306468
rect 299532 306428 300032 306456
rect 299532 306416 299538 306428
rect 300026 306416 300032 306428
rect 300084 306416 300090 306468
rect 302234 306416 302240 306468
rect 302292 306456 302298 306468
rect 302694 306456 302700 306468
rect 302292 306428 302700 306456
rect 302292 306416 302298 306428
rect 302694 306416 302700 306428
rect 302752 306416 302758 306468
rect 306466 306416 306472 306468
rect 306524 306456 306530 306468
rect 306742 306456 306748 306468
rect 306524 306428 306748 306456
rect 306524 306416 306530 306428
rect 306742 306416 306748 306428
rect 306800 306416 306806 306468
rect 312262 306416 312268 306468
rect 312320 306456 312326 306468
rect 312630 306456 312636 306468
rect 312320 306428 312636 306456
rect 312320 306416 312326 306428
rect 312630 306416 312636 306428
rect 312688 306416 312694 306468
rect 313274 306416 313280 306468
rect 313332 306456 313338 306468
rect 314194 306456 314200 306468
rect 313332 306428 314200 306456
rect 313332 306416 313338 306428
rect 314194 306416 314200 306428
rect 314252 306416 314258 306468
rect 316034 306416 316040 306468
rect 316092 306456 316098 306468
rect 316770 306456 316776 306468
rect 316092 306428 316776 306456
rect 316092 306416 316098 306428
rect 316770 306416 316776 306428
rect 316828 306416 316834 306468
rect 322934 306416 322940 306468
rect 322992 306456 322998 306468
rect 323486 306456 323492 306468
rect 322992 306428 323492 306456
rect 322992 306416 322998 306428
rect 323486 306416 323492 306428
rect 323544 306416 323550 306468
rect 325694 306416 325700 306468
rect 325752 306456 325758 306468
rect 326154 306456 326160 306468
rect 325752 306428 326160 306456
rect 325752 306416 325758 306428
rect 326154 306416 326160 306428
rect 326212 306416 326218 306468
rect 327074 306416 327080 306468
rect 327132 306456 327138 306468
rect 327902 306456 327908 306468
rect 327132 306428 327908 306456
rect 327132 306416 327138 306428
rect 327902 306416 327908 306428
rect 327960 306416 327966 306468
rect 329834 306416 329840 306468
rect 329892 306456 329898 306468
rect 330662 306456 330668 306468
rect 329892 306428 330668 306456
rect 329892 306416 329898 306428
rect 330662 306416 330668 306428
rect 330720 306416 330726 306468
rect 331950 306456 331956 306468
rect 331232 306428 331956 306456
rect 241790 306348 241796 306400
rect 241848 306388 241854 306400
rect 242526 306388 242532 306400
rect 241848 306360 242532 306388
rect 241848 306348 241854 306360
rect 242526 306348 242532 306360
rect 242584 306348 242590 306400
rect 247402 306348 247408 306400
rect 247460 306388 247466 306400
rect 248322 306388 248328 306400
rect 247460 306360 248328 306388
rect 247460 306348 247466 306360
rect 248322 306348 248328 306360
rect 248380 306348 248386 306400
rect 248506 306348 248512 306400
rect 248564 306388 248570 306400
rect 249242 306388 249248 306400
rect 248564 306360 249248 306388
rect 248564 306348 248570 306360
rect 249242 306348 249248 306360
rect 249300 306348 249306 306400
rect 259546 306348 259552 306400
rect 259604 306388 259610 306400
rect 260558 306388 260564 306400
rect 259604 306360 260564 306388
rect 259604 306348 259610 306360
rect 260558 306348 260564 306360
rect 260616 306348 260622 306400
rect 262398 306348 262404 306400
rect 262456 306388 262462 306400
rect 262950 306388 262956 306400
rect 262456 306360 262956 306388
rect 262456 306348 262462 306360
rect 262950 306348 262956 306360
rect 263008 306348 263014 306400
rect 266814 306348 266820 306400
rect 266872 306388 266878 306400
rect 267458 306388 267464 306400
rect 266872 306360 267464 306388
rect 266872 306348 266878 306360
rect 267458 306348 267464 306360
rect 267516 306348 267522 306400
rect 267734 306348 267740 306400
rect 267792 306388 267798 306400
rect 268378 306388 268384 306400
rect 267792 306360 268384 306388
rect 267792 306348 267798 306360
rect 268378 306348 268384 306360
rect 268436 306348 268442 306400
rect 269390 306348 269396 306400
rect 269448 306388 269454 306400
rect 270034 306388 270040 306400
rect 269448 306360 270040 306388
rect 269448 306348 269454 306360
rect 270034 306348 270040 306360
rect 270092 306348 270098 306400
rect 272150 306348 272156 306400
rect 272208 306388 272214 306400
rect 272518 306388 272524 306400
rect 272208 306360 272524 306388
rect 272208 306348 272214 306360
rect 272518 306348 272524 306360
rect 272576 306348 272582 306400
rect 285766 306348 285772 306400
rect 285824 306388 285830 306400
rect 286134 306388 286140 306400
rect 285824 306360 286140 306388
rect 285824 306348 285830 306360
rect 286134 306348 286140 306360
rect 286192 306348 286198 306400
rect 287422 306348 287428 306400
rect 287480 306388 287486 306400
rect 288158 306388 288164 306400
rect 287480 306360 288164 306388
rect 287480 306348 287486 306360
rect 288158 306348 288164 306360
rect 288216 306348 288222 306400
rect 288434 306348 288440 306400
rect 288492 306388 288498 306400
rect 289262 306388 289268 306400
rect 288492 306360 289268 306388
rect 288492 306348 288498 306360
rect 289262 306348 289268 306360
rect 289320 306348 289326 306400
rect 289814 306348 289820 306400
rect 289872 306388 289878 306400
rect 290090 306388 290096 306400
rect 289872 306360 290096 306388
rect 289872 306348 289878 306360
rect 290090 306348 290096 306360
rect 290148 306348 290154 306400
rect 291194 306348 291200 306400
rect 291252 306388 291258 306400
rect 291562 306388 291568 306400
rect 291252 306360 291568 306388
rect 291252 306348 291258 306360
rect 291562 306348 291568 306360
rect 291620 306348 291626 306400
rect 291654 306348 291660 306400
rect 291712 306388 291718 306400
rect 292206 306388 292212 306400
rect 291712 306360 292212 306388
rect 291712 306348 291718 306360
rect 292206 306348 292212 306360
rect 292264 306348 292270 306400
rect 292850 306348 292856 306400
rect 292908 306388 292914 306400
rect 293402 306388 293408 306400
rect 292908 306360 293408 306388
rect 292908 306348 292914 306360
rect 293402 306348 293408 306360
rect 293460 306348 293466 306400
rect 294138 306348 294144 306400
rect 294196 306388 294202 306400
rect 294598 306388 294604 306400
rect 294196 306360 294604 306388
rect 294196 306348 294202 306360
rect 294598 306348 294604 306360
rect 294656 306348 294662 306400
rect 295518 306348 295524 306400
rect 295576 306388 295582 306400
rect 295978 306388 295984 306400
rect 295576 306360 295984 306388
rect 295576 306348 295582 306360
rect 295978 306348 295984 306360
rect 296036 306348 296042 306400
rect 296714 306348 296720 306400
rect 296772 306388 296778 306400
rect 297450 306388 297456 306400
rect 296772 306360 297456 306388
rect 296772 306348 296778 306360
rect 297450 306348 297456 306360
rect 297508 306348 297514 306400
rect 298094 306348 298100 306400
rect 298152 306388 298158 306400
rect 298554 306388 298560 306400
rect 298152 306360 298560 306388
rect 298152 306348 298158 306360
rect 298554 306348 298560 306360
rect 298612 306348 298618 306400
rect 299750 306348 299756 306400
rect 299808 306388 299814 306400
rect 300578 306388 300584 306400
rect 299808 306360 300584 306388
rect 299808 306348 299814 306360
rect 300578 306348 300584 306360
rect 300636 306348 300642 306400
rect 301222 306348 301228 306400
rect 301280 306388 301286 306400
rect 301774 306388 301780 306400
rect 301280 306360 301780 306388
rect 301280 306348 301286 306360
rect 301774 306348 301780 306360
rect 301832 306348 301838 306400
rect 302510 306348 302516 306400
rect 302568 306388 302574 306400
rect 302878 306388 302884 306400
rect 302568 306360 302884 306388
rect 302568 306348 302574 306360
rect 302878 306348 302884 306360
rect 302936 306348 302942 306400
rect 303706 306348 303712 306400
rect 303764 306388 303770 306400
rect 304626 306388 304632 306400
rect 303764 306360 304632 306388
rect 303764 306348 303770 306360
rect 304626 306348 304632 306360
rect 304684 306348 304690 306400
rect 306558 306348 306564 306400
rect 306616 306388 306622 306400
rect 307202 306388 307208 306400
rect 306616 306360 307208 306388
rect 306616 306348 306622 306360
rect 307202 306348 307208 306360
rect 307260 306348 307266 306400
rect 307754 306348 307760 306400
rect 307812 306388 307818 306400
rect 308398 306388 308404 306400
rect 307812 306360 308404 306388
rect 307812 306348 307818 306360
rect 308398 306348 308404 306360
rect 308456 306348 308462 306400
rect 309134 306348 309140 306400
rect 309192 306388 309198 306400
rect 310054 306388 310060 306400
rect 309192 306360 310060 306388
rect 309192 306348 309198 306360
rect 310054 306348 310060 306360
rect 310112 306348 310118 306400
rect 310698 306348 310704 306400
rect 310756 306388 310762 306400
rect 311802 306388 311808 306400
rect 310756 306360 311808 306388
rect 310756 306348 310762 306360
rect 311802 306348 311808 306360
rect 311860 306348 311866 306400
rect 313458 306348 313464 306400
rect 313516 306388 313522 306400
rect 314378 306388 314384 306400
rect 313516 306360 314384 306388
rect 313516 306348 313522 306360
rect 314378 306348 314384 306360
rect 314436 306348 314442 306400
rect 314838 306348 314844 306400
rect 314896 306388 314902 306400
rect 315298 306388 315304 306400
rect 314896 306360 315304 306388
rect 314896 306348 314902 306360
rect 315298 306348 315304 306360
rect 315356 306348 315362 306400
rect 316218 306348 316224 306400
rect 316276 306388 316282 306400
rect 316862 306388 316868 306400
rect 316276 306360 316868 306388
rect 316276 306348 316282 306360
rect 316862 306348 316868 306360
rect 316920 306348 316926 306400
rect 317414 306348 317420 306400
rect 317472 306388 317478 306400
rect 317966 306388 317972 306400
rect 317472 306360 317972 306388
rect 317472 306348 317478 306360
rect 317966 306348 317972 306360
rect 318024 306348 318030 306400
rect 318886 306348 318892 306400
rect 318944 306388 318950 306400
rect 319806 306388 319812 306400
rect 318944 306360 319812 306388
rect 318944 306348 318950 306360
rect 319806 306348 319812 306360
rect 319864 306348 319870 306400
rect 320450 306348 320456 306400
rect 320508 306388 320514 306400
rect 321370 306388 321376 306400
rect 320508 306360 321376 306388
rect 320508 306348 320514 306360
rect 321370 306348 321376 306360
rect 321428 306348 321434 306400
rect 324314 306348 324320 306400
rect 324372 306388 324378 306400
rect 325050 306388 325056 306400
rect 324372 306360 325056 306388
rect 324372 306348 324378 306360
rect 325050 306348 325056 306360
rect 325108 306348 325114 306400
rect 325878 306348 325884 306400
rect 325936 306388 325942 306400
rect 326430 306388 326436 306400
rect 325936 306360 326436 306388
rect 325936 306348 325942 306360
rect 326430 306348 326436 306360
rect 326488 306348 326494 306400
rect 327442 306348 327448 306400
rect 327500 306388 327506 306400
rect 328086 306388 328092 306400
rect 327500 306360 328092 306388
rect 327500 306348 327506 306360
rect 328086 306348 328092 306360
rect 328144 306348 328150 306400
rect 328454 306348 328460 306400
rect 328512 306388 328518 306400
rect 329190 306388 329196 306400
rect 328512 306360 329196 306388
rect 328512 306348 328518 306360
rect 329190 306348 329196 306360
rect 329248 306348 329254 306400
rect 241698 306280 241704 306332
rect 241756 306320 241762 306332
rect 242434 306320 242440 306332
rect 241756 306292 242440 306320
rect 241756 306280 241762 306292
rect 242434 306280 242440 306292
rect 242492 306280 242498 306332
rect 247310 306280 247316 306332
rect 247368 306320 247374 306332
rect 247862 306320 247868 306332
rect 247368 306292 247868 306320
rect 247368 306280 247374 306292
rect 247862 306280 247868 306292
rect 247920 306280 247926 306332
rect 248690 306280 248696 306332
rect 248748 306320 248754 306332
rect 249150 306320 249156 306332
rect 248748 306292 249156 306320
rect 248748 306280 248754 306292
rect 249150 306280 249156 306292
rect 249208 306280 249214 306332
rect 249886 306280 249892 306332
rect 249944 306320 249950 306332
rect 250714 306320 250720 306332
rect 249944 306292 250720 306320
rect 249944 306280 249950 306292
rect 250714 306280 250720 306292
rect 250772 306280 250778 306332
rect 252738 306280 252744 306332
rect 252796 306320 252802 306332
rect 253750 306320 253756 306332
rect 252796 306292 253756 306320
rect 252796 306280 252802 306292
rect 253750 306280 253756 306292
rect 253808 306280 253814 306332
rect 254210 306280 254216 306332
rect 254268 306320 254274 306332
rect 255038 306320 255044 306332
rect 254268 306292 255044 306320
rect 254268 306280 254274 306292
rect 255038 306280 255044 306292
rect 255096 306280 255102 306332
rect 255774 306280 255780 306332
rect 255832 306320 255838 306332
rect 256326 306320 256332 306332
rect 255832 306292 256332 306320
rect 255832 306280 255838 306292
rect 256326 306280 256332 306292
rect 256384 306280 256390 306332
rect 256878 306280 256884 306332
rect 256936 306320 256942 306332
rect 257430 306320 257436 306332
rect 256936 306292 257436 306320
rect 256936 306280 256942 306292
rect 257430 306280 257436 306292
rect 257488 306280 257494 306332
rect 258166 306280 258172 306332
rect 258224 306320 258230 306332
rect 259178 306320 259184 306332
rect 258224 306292 259184 306320
rect 258224 306280 258230 306292
rect 259178 306280 259184 306292
rect 259236 306280 259242 306332
rect 259730 306280 259736 306332
rect 259788 306320 259794 306332
rect 260466 306320 260472 306332
rect 259788 306292 260472 306320
rect 259788 306280 259794 306292
rect 260466 306280 260472 306292
rect 260524 306280 260530 306332
rect 262582 306280 262588 306332
rect 262640 306320 262646 306332
rect 263502 306320 263508 306332
rect 262640 306292 263508 306320
rect 262640 306280 262646 306292
rect 263502 306280 263508 306292
rect 263560 306280 263566 306332
rect 263686 306280 263692 306332
rect 263744 306320 263750 306332
rect 263962 306320 263968 306332
rect 263744 306292 263968 306320
rect 263744 306280 263750 306292
rect 263962 306280 263968 306292
rect 264020 306280 264026 306332
rect 265342 306280 265348 306332
rect 265400 306320 265406 306332
rect 265986 306320 265992 306332
rect 265400 306292 265992 306320
rect 265400 306280 265406 306292
rect 265986 306280 265992 306292
rect 266044 306280 266050 306332
rect 266630 306280 266636 306332
rect 266688 306320 266694 306332
rect 266998 306320 267004 306332
rect 266688 306292 267004 306320
rect 266688 306280 266694 306292
rect 266998 306280 267004 306292
rect 267056 306280 267062 306332
rect 268010 306280 268016 306332
rect 268068 306320 268074 306332
rect 268838 306320 268844 306332
rect 268068 306292 268844 306320
rect 268068 306280 268074 306292
rect 268838 306280 268844 306292
rect 268896 306280 268902 306332
rect 269298 306280 269304 306332
rect 269356 306320 269362 306332
rect 269850 306320 269856 306332
rect 269356 306292 269856 306320
rect 269356 306280 269362 306292
rect 269850 306280 269856 306292
rect 269908 306280 269914 306332
rect 271966 306280 271972 306332
rect 272024 306320 272030 306332
rect 272426 306320 272432 306332
rect 272024 306292 272432 306320
rect 272024 306280 272030 306292
rect 272426 306280 272432 306292
rect 272484 306280 272490 306332
rect 273254 306280 273260 306332
rect 273312 306320 273318 306332
rect 274174 306320 274180 306332
rect 273312 306292 274180 306320
rect 273312 306280 273318 306292
rect 274174 306280 274180 306292
rect 274232 306280 274238 306332
rect 274726 306280 274732 306332
rect 274784 306320 274790 306332
rect 274910 306320 274916 306332
rect 274784 306292 274916 306320
rect 274784 306280 274790 306292
rect 274910 306280 274916 306292
rect 274968 306280 274974 306332
rect 277394 306280 277400 306332
rect 277452 306320 277458 306332
rect 278498 306320 278504 306332
rect 277452 306292 278504 306320
rect 277452 306280 277458 306292
rect 278498 306280 278504 306292
rect 278556 306280 278562 306332
rect 280430 306280 280436 306332
rect 280488 306320 280494 306332
rect 280890 306320 280896 306332
rect 280488 306292 280896 306320
rect 280488 306280 280494 306292
rect 280890 306280 280896 306292
rect 280948 306280 280954 306332
rect 280982 306280 280988 306332
rect 281040 306320 281046 306332
rect 331232 306320 331260 306428
rect 331950 306416 331956 306428
rect 332008 306416 332014 306468
rect 332686 306416 332692 306468
rect 332744 306456 332750 306468
rect 333054 306456 333060 306468
rect 332744 306428 333060 306456
rect 332744 306416 332750 306428
rect 333054 306416 333060 306428
rect 333112 306416 333118 306468
rect 333974 306348 333980 306400
rect 334032 306388 334038 306400
rect 335078 306388 335084 306400
rect 334032 306360 335084 306388
rect 334032 306348 334038 306360
rect 335078 306348 335084 306360
rect 335136 306348 335142 306400
rect 335630 306348 335636 306400
rect 335688 306388 335694 306400
rect 336550 306388 336556 306400
rect 335688 306360 336556 306388
rect 335688 306348 335694 306360
rect 336550 306348 336556 306360
rect 336608 306348 336614 306400
rect 281040 306292 331260 306320
rect 281040 306280 281046 306292
rect 331306 306280 331312 306332
rect 331364 306320 331370 306332
rect 332318 306320 332324 306332
rect 331364 306292 332324 306320
rect 331364 306280 331370 306292
rect 332318 306280 332324 306292
rect 332376 306280 332382 306332
rect 332594 306280 332600 306332
rect 332652 306320 332658 306332
rect 333606 306320 333612 306332
rect 332652 306292 333612 306320
rect 332652 306280 332658 306292
rect 333606 306280 333612 306292
rect 333664 306280 333670 306332
rect 334066 306280 334072 306332
rect 334124 306320 334130 306332
rect 334710 306320 334716 306332
rect 334124 306292 334716 306320
rect 334124 306280 334130 306292
rect 334710 306280 334716 306292
rect 334768 306280 334774 306332
rect 335722 306280 335728 306332
rect 335780 306320 335786 306332
rect 335998 306320 336004 306332
rect 335780 306292 336004 306320
rect 335780 306280 335786 306292
rect 335998 306280 336004 306292
rect 336056 306280 336062 306332
rect 336918 306280 336924 306332
rect 336976 306320 336982 306332
rect 337102 306320 337108 306332
rect 336976 306292 337108 306320
rect 336976 306280 336982 306292
rect 337102 306280 337108 306292
rect 337160 306280 337166 306332
rect 338206 306280 338212 306332
rect 338264 306320 338270 306332
rect 339402 306320 339408 306332
rect 338264 306292 339408 306320
rect 338264 306280 338270 306292
rect 339402 306280 339408 306292
rect 339460 306280 339466 306332
rect 339586 306280 339592 306332
rect 339644 306320 339650 306332
rect 340690 306320 340696 306332
rect 339644 306292 340696 306320
rect 339644 306280 339650 306292
rect 340690 306280 340696 306292
rect 340748 306280 340754 306332
rect 230934 306212 230940 306264
rect 230992 306252 230998 306264
rect 231578 306252 231584 306264
rect 230992 306224 231584 306252
rect 230992 306212 230998 306224
rect 231578 306212 231584 306224
rect 231636 306212 231642 306264
rect 237466 306212 237472 306264
rect 237524 306252 237530 306264
rect 237926 306252 237932 306264
rect 237524 306224 237932 306252
rect 237524 306212 237530 306224
rect 237926 306212 237932 306224
rect 237984 306212 237990 306264
rect 238846 306212 238852 306264
rect 238904 306212 238910 306264
rect 239030 306212 239036 306264
rect 239088 306252 239094 306264
rect 239674 306252 239680 306264
rect 239088 306224 239680 306252
rect 239088 306212 239094 306224
rect 239674 306212 239680 306224
rect 239732 306212 239738 306264
rect 240410 306212 240416 306264
rect 240468 306252 240474 306264
rect 241330 306252 241336 306264
rect 240468 306224 241336 306252
rect 240468 306212 240474 306224
rect 241330 306212 241336 306224
rect 241388 306212 241394 306264
rect 243170 306212 243176 306264
rect 243228 306252 243234 306264
rect 244182 306252 244188 306264
rect 243228 306224 244188 306252
rect 243228 306212 243234 306224
rect 244182 306212 244188 306224
rect 244240 306212 244246 306264
rect 244734 306212 244740 306264
rect 244792 306252 244798 306264
rect 245470 306252 245476 306264
rect 244792 306224 245476 306252
rect 244792 306212 244798 306224
rect 245470 306212 245476 306224
rect 245528 306212 245534 306264
rect 246022 306212 246028 306264
rect 246080 306252 246086 306264
rect 246758 306252 246764 306264
rect 246080 306224 246764 306252
rect 246080 306212 246086 306224
rect 246758 306212 246764 306224
rect 246816 306212 246822 306264
rect 247494 306212 247500 306264
rect 247552 306252 247558 306264
rect 247954 306252 247960 306264
rect 247552 306224 247960 306252
rect 247552 306212 247558 306224
rect 247954 306212 247960 306224
rect 248012 306212 248018 306264
rect 250070 306212 250076 306264
rect 250128 306252 250134 306264
rect 250898 306252 250904 306264
rect 250128 306224 250904 306252
rect 250128 306212 250134 306224
rect 250898 306212 250904 306224
rect 250956 306212 250962 306264
rect 262306 306212 262312 306264
rect 262364 306252 262370 306264
rect 263318 306252 263324 306264
rect 262364 306224 263324 306252
rect 262364 306212 262370 306224
rect 263318 306212 263324 306224
rect 263376 306212 263382 306264
rect 265250 306212 265256 306264
rect 265308 306252 265314 306264
rect 265710 306252 265716 306264
rect 265308 306224 265716 306252
rect 265308 306212 265314 306224
rect 265710 306212 265716 306224
rect 265768 306212 265774 306264
rect 266538 306212 266544 306264
rect 266596 306252 266602 306264
rect 267642 306252 267648 306264
rect 266596 306224 267648 306252
rect 266596 306212 266602 306224
rect 267642 306212 267648 306224
rect 267700 306212 267706 306264
rect 268102 306212 268108 306264
rect 268160 306252 268166 306264
rect 268746 306252 268752 306264
rect 268160 306224 268752 306252
rect 268160 306212 268166 306224
rect 268746 306212 268752 306224
rect 268804 306212 268810 306264
rect 269206 306212 269212 306264
rect 269264 306252 269270 306264
rect 270126 306252 270132 306264
rect 269264 306224 270132 306252
rect 269264 306212 269270 306224
rect 270126 306212 270132 306224
rect 270184 306212 270190 306264
rect 270678 306212 270684 306264
rect 270736 306252 270742 306264
rect 271046 306252 271052 306264
rect 270736 306224 271052 306252
rect 270736 306212 270742 306224
rect 271046 306212 271052 306224
rect 271104 306212 271110 306264
rect 273346 306212 273352 306264
rect 273404 306252 273410 306264
rect 273714 306252 273720 306264
rect 273404 306224 273720 306252
rect 273404 306212 273410 306224
rect 273714 306212 273720 306224
rect 273772 306212 273778 306264
rect 277578 306212 277584 306264
rect 277636 306252 277642 306264
rect 278314 306252 278320 306264
rect 277636 306224 278320 306252
rect 277636 306212 277642 306224
rect 278314 306212 278320 306224
rect 278372 306212 278378 306264
rect 340966 306252 340972 306264
rect 279988 306224 340972 306252
rect 237742 306144 237748 306196
rect 237800 306184 237806 306196
rect 238386 306184 238392 306196
rect 237800 306156 238392 306184
rect 237800 306144 237806 306156
rect 238386 306144 238392 306156
rect 238444 306144 238450 306196
rect 238754 306144 238760 306196
rect 238812 306184 238818 306196
rect 240042 306184 240048 306196
rect 238812 306156 240048 306184
rect 238812 306144 238818 306156
rect 240042 306144 240048 306156
rect 240100 306144 240106 306196
rect 257062 306144 257068 306196
rect 257120 306184 257126 306196
rect 257522 306184 257528 306196
rect 257120 306156 257528 306184
rect 257120 306144 257126 306156
rect 257522 306144 257528 306156
rect 257580 306144 257586 306196
rect 258350 306144 258356 306196
rect 258408 306184 258414 306196
rect 258810 306184 258816 306196
rect 258408 306156 258816 306184
rect 258408 306144 258414 306156
rect 258810 306144 258816 306156
rect 258868 306144 258874 306196
rect 259454 306144 259460 306196
rect 259512 306184 259518 306196
rect 260006 306184 260012 306196
rect 259512 306156 260012 306184
rect 259512 306144 259518 306156
rect 260006 306144 260012 306156
rect 260064 306144 260070 306196
rect 270862 306144 270868 306196
rect 270920 306144 270926 306196
rect 274910 306144 274916 306196
rect 274968 306184 274974 306196
rect 275922 306184 275928 306196
rect 274968 306156 275928 306184
rect 274968 306144 274974 306156
rect 275922 306144 275928 306156
rect 275980 306144 275986 306196
rect 276934 306144 276940 306196
rect 276992 306184 276998 306196
rect 279988 306184 280016 306224
rect 340966 306212 340972 306224
rect 341024 306212 341030 306264
rect 342254 306184 342260 306196
rect 276992 306156 280016 306184
rect 280080 306156 342260 306184
rect 276992 306144 276998 306156
rect 237558 306076 237564 306128
rect 237616 306116 237622 306128
rect 238294 306116 238300 306128
rect 237616 306088 238300 306116
rect 237616 306076 237622 306088
rect 238294 306076 238300 306088
rect 238352 306076 238358 306128
rect 255498 306076 255504 306128
rect 255556 306116 255562 306128
rect 255958 306116 255964 306128
rect 255556 306088 255964 306116
rect 255556 306076 255562 306088
rect 255958 306076 255964 306088
rect 256016 306076 256022 306128
rect 256786 306076 256792 306128
rect 256844 306116 256850 306128
rect 257890 306116 257896 306128
rect 256844 306088 257896 306116
rect 256844 306076 256850 306088
rect 257890 306076 257896 306088
rect 257948 306076 257954 306128
rect 263962 306076 263968 306128
rect 264020 306116 264026 306128
rect 264698 306116 264704 306128
rect 264020 306088 264704 306116
rect 264020 306076 264026 306088
rect 264698 306076 264704 306088
rect 264756 306076 264762 306128
rect 255406 306008 255412 306060
rect 255464 306048 255470 306060
rect 256418 306048 256424 306060
rect 255464 306020 256424 306048
rect 255464 306008 255470 306020
rect 256418 306008 256424 306020
rect 256476 306008 256482 306060
rect 230842 305940 230848 305992
rect 230900 305980 230906 305992
rect 231118 305980 231124 305992
rect 230900 305952 231124 305980
rect 230900 305940 230906 305952
rect 231118 305940 231124 305952
rect 231176 305940 231182 305992
rect 263778 305940 263784 305992
rect 263836 305980 263842 305992
rect 264422 305980 264428 305992
rect 263836 305952 264428 305980
rect 263836 305940 263842 305952
rect 264422 305940 264428 305952
rect 264480 305940 264486 305992
rect 270586 305940 270592 305992
rect 270644 305980 270650 305992
rect 270880 305980 270908 306144
rect 277026 306076 277032 306128
rect 277084 306116 277090 306128
rect 280080 306116 280108 306156
rect 342254 306144 342260 306156
rect 342312 306144 342318 306196
rect 280982 306116 280988 306128
rect 277084 306088 280108 306116
rect 280172 306088 280988 306116
rect 277084 306076 277090 306088
rect 277118 306008 277124 306060
rect 277176 306048 277182 306060
rect 280172 306048 280200 306088
rect 280982 306076 280988 306088
rect 281040 306076 281046 306128
rect 281718 306076 281724 306128
rect 281776 306116 281782 306128
rect 282454 306116 282460 306128
rect 281776 306088 282460 306116
rect 281776 306076 281782 306088
rect 282454 306076 282460 306088
rect 282512 306076 282518 306128
rect 282730 306076 282736 306128
rect 282788 306116 282794 306128
rect 350626 306116 350632 306128
rect 282788 306088 350632 306116
rect 282788 306076 282794 306088
rect 350626 306076 350632 306088
rect 350684 306076 350690 306128
rect 277176 306020 280200 306048
rect 277176 306008 277182 306020
rect 282638 306008 282644 306060
rect 282696 306048 282702 306060
rect 354858 306048 354864 306060
rect 282696 306020 354864 306048
rect 282696 306008 282702 306020
rect 354858 306008 354864 306020
rect 354916 306008 354922 306060
rect 270644 305952 270908 305980
rect 270644 305940 270650 305952
rect 281074 305940 281080 305992
rect 281132 305980 281138 305992
rect 354214 305980 354220 305992
rect 281132 305952 354220 305980
rect 281132 305940 281138 305952
rect 354214 305940 354220 305952
rect 354272 305940 354278 305992
rect 270678 305872 270684 305924
rect 270736 305912 270742 305924
rect 271598 305912 271604 305924
rect 270736 305884 271604 305912
rect 270736 305872 270742 305884
rect 271598 305872 271604 305884
rect 271656 305872 271662 305924
rect 280982 305872 280988 305924
rect 281040 305912 281046 305924
rect 354674 305912 354680 305924
rect 281040 305884 354680 305912
rect 281040 305872 281046 305884
rect 354674 305872 354680 305884
rect 354732 305872 354738 305924
rect 270494 305804 270500 305856
rect 270552 305844 270558 305856
rect 271782 305844 271788 305856
rect 270552 305816 271788 305844
rect 270552 305804 270558 305816
rect 271782 305804 271788 305816
rect 271840 305804 271846 305856
rect 280890 305804 280896 305856
rect 280948 305844 280954 305856
rect 354766 305844 354772 305856
rect 280948 305816 354772 305844
rect 280948 305804 280954 305816
rect 354766 305804 354772 305816
rect 354824 305804 354830 305856
rect 280798 305736 280804 305788
rect 280856 305776 280862 305788
rect 356146 305776 356152 305788
rect 280856 305748 356152 305776
rect 280856 305736 280862 305748
rect 356146 305736 356152 305748
rect 356204 305736 356210 305788
rect 75914 305668 75920 305720
rect 75972 305708 75978 305720
rect 243998 305708 244004 305720
rect 75972 305680 244004 305708
rect 75972 305668 75978 305680
rect 243998 305668 244004 305680
rect 244056 305668 244062 305720
rect 277302 305668 277308 305720
rect 277360 305708 277366 305720
rect 353662 305708 353668 305720
rect 277360 305680 353668 305708
rect 277360 305668 277366 305680
rect 353662 305668 353668 305680
rect 353720 305668 353726 305720
rect 72418 305600 72424 305652
rect 72476 305640 72482 305652
rect 242986 305640 242992 305652
rect 72476 305612 242992 305640
rect 72476 305600 72482 305612
rect 242986 305600 242992 305612
rect 243044 305600 243050 305652
rect 278314 305600 278320 305652
rect 278372 305640 278378 305652
rect 357434 305640 357440 305652
rect 278372 305612 357440 305640
rect 278372 305600 278378 305612
rect 357434 305600 357440 305612
rect 357492 305600 357498 305652
rect 283006 305532 283012 305584
rect 283064 305572 283070 305584
rect 284202 305572 284208 305584
rect 283064 305544 284208 305572
rect 283064 305532 283070 305544
rect 284202 305532 284208 305544
rect 284260 305532 284266 305584
rect 284386 305532 284392 305584
rect 284444 305572 284450 305584
rect 285122 305572 285128 305584
rect 284444 305544 285128 305572
rect 284444 305532 284450 305544
rect 285122 305532 285128 305544
rect 285180 305532 285186 305584
rect 287238 305532 287244 305584
rect 287296 305572 287302 305584
rect 287882 305572 287888 305584
rect 287296 305544 287888 305572
rect 287296 305532 287302 305544
rect 287882 305532 287888 305544
rect 287940 305532 287946 305584
rect 288618 305532 288624 305584
rect 288676 305572 288682 305584
rect 289170 305572 289176 305584
rect 288676 305544 289176 305572
rect 288676 305532 288682 305544
rect 289170 305532 289176 305544
rect 289228 305532 289234 305584
rect 289998 305532 290004 305584
rect 290056 305572 290062 305584
rect 290458 305572 290464 305584
rect 290056 305544 290464 305572
rect 290056 305532 290062 305544
rect 290458 305532 290464 305544
rect 290516 305532 290522 305584
rect 291194 305532 291200 305584
rect 291252 305572 291258 305584
rect 292022 305572 292028 305584
rect 291252 305544 292028 305572
rect 291252 305532 291258 305544
rect 292022 305532 292028 305544
rect 292080 305532 292086 305584
rect 332502 305572 332508 305584
rect 292546 305544 332508 305572
rect 284478 305464 284484 305516
rect 284536 305504 284542 305516
rect 285030 305504 285036 305516
rect 284536 305476 285036 305504
rect 284536 305464 284542 305476
rect 285030 305464 285036 305476
rect 285088 305464 285094 305516
rect 287054 305464 287060 305516
rect 287112 305504 287118 305516
rect 288066 305504 288072 305516
rect 287112 305476 288072 305504
rect 287112 305464 287118 305476
rect 288066 305464 288072 305476
rect 288124 305464 288130 305516
rect 288802 305464 288808 305516
rect 288860 305504 288866 305516
rect 289630 305504 289636 305516
rect 288860 305476 289636 305504
rect 288860 305464 288866 305476
rect 289630 305464 289636 305476
rect 289688 305464 289694 305516
rect 289814 305464 289820 305516
rect 289872 305504 289878 305516
rect 290550 305504 290556 305516
rect 289872 305476 290556 305504
rect 289872 305464 289878 305476
rect 290550 305464 290556 305476
rect 290608 305464 290614 305516
rect 283926 305396 283932 305448
rect 283984 305436 283990 305448
rect 284202 305436 284208 305448
rect 283984 305408 284208 305436
rect 283984 305396 283990 305408
rect 284202 305396 284208 305408
rect 284260 305396 284266 305448
rect 289538 305396 289544 305448
rect 289596 305436 289602 305448
rect 292546 305436 292574 305544
rect 332502 305532 332508 305544
rect 332560 305532 332566 305584
rect 332870 305532 332876 305584
rect 332928 305572 332934 305584
rect 333330 305572 333336 305584
rect 332928 305544 333336 305572
rect 332928 305532 332934 305544
rect 333330 305532 333336 305544
rect 333388 305532 333394 305584
rect 334250 305532 334256 305584
rect 334308 305572 334314 305584
rect 335262 305572 335268 305584
rect 334308 305544 335268 305572
rect 334308 305532 334314 305544
rect 335262 305532 335268 305544
rect 335320 305532 335326 305584
rect 335538 305532 335544 305584
rect 335596 305572 335602 305584
rect 336366 305572 336372 305584
rect 335596 305544 336372 305572
rect 335596 305532 335602 305544
rect 336366 305532 336372 305544
rect 336424 305532 336430 305584
rect 339678 305532 339684 305584
rect 339736 305572 339742 305584
rect 340138 305572 340144 305584
rect 339736 305544 340144 305572
rect 339736 305532 339742 305544
rect 340138 305532 340144 305544
rect 340196 305532 340202 305584
rect 294230 305464 294236 305516
rect 294288 305504 294294 305516
rect 294690 305504 294696 305516
rect 294288 305476 294696 305504
rect 294288 305464 294294 305476
rect 294690 305464 294696 305476
rect 294748 305464 294754 305516
rect 295794 305464 295800 305516
rect 295852 305504 295858 305516
rect 295978 305504 295984 305516
rect 295852 305476 295984 305504
rect 295852 305464 295858 305476
rect 295978 305464 295984 305476
rect 296036 305464 296042 305516
rect 299842 305464 299848 305516
rect 299900 305504 299906 305516
rect 300486 305504 300492 305516
rect 299900 305476 300492 305504
rect 299900 305464 299906 305476
rect 300486 305464 300492 305476
rect 300544 305464 300550 305516
rect 300946 305464 300952 305516
rect 301004 305504 301010 305516
rect 301590 305504 301596 305516
rect 301004 305476 301596 305504
rect 301004 305464 301010 305476
rect 301590 305464 301596 305476
rect 301648 305464 301654 305516
rect 340874 305504 340880 305516
rect 301976 305476 331444 305504
rect 289596 305408 292574 305436
rect 289596 305396 289602 305408
rect 301038 305396 301044 305448
rect 301096 305436 301102 305448
rect 301866 305436 301872 305448
rect 301096 305408 301872 305436
rect 301096 305396 301102 305408
rect 301866 305396 301872 305408
rect 301924 305396 301930 305448
rect 236638 305328 236644 305380
rect 236696 305368 236702 305380
rect 236822 305368 236828 305380
rect 236696 305340 236828 305368
rect 236696 305328 236702 305340
rect 236822 305328 236828 305340
rect 236880 305328 236886 305380
rect 295058 305260 295064 305312
rect 295116 305300 295122 305312
rect 301976 305300 302004 305476
rect 331416 305436 331444 305476
rect 331600 305476 340880 305504
rect 331600 305436 331628 305476
rect 340874 305464 340880 305476
rect 340932 305464 340938 305516
rect 295116 305272 302004 305300
rect 302206 305408 331260 305436
rect 331416 305408 331628 305436
rect 295116 305260 295122 305272
rect 260926 305192 260932 305244
rect 260984 305232 260990 305244
rect 262030 305232 262036 305244
rect 260984 305204 262036 305232
rect 260984 305192 260990 305204
rect 262030 305192 262036 305204
rect 262088 305192 262094 305244
rect 298002 305192 298008 305244
rect 298060 305232 298066 305244
rect 302206 305232 302234 305408
rect 303798 305328 303804 305380
rect 303856 305368 303862 305380
rect 304810 305368 304816 305380
rect 303856 305340 304816 305368
rect 303856 305328 303862 305340
rect 304810 305328 304816 305340
rect 304868 305328 304874 305380
rect 305270 305328 305276 305380
rect 305328 305368 305334 305380
rect 306006 305368 306012 305380
rect 305328 305340 306012 305368
rect 305328 305328 305334 305340
rect 306006 305328 306012 305340
rect 306064 305328 306070 305380
rect 306374 305328 306380 305380
rect 306432 305368 306438 305380
rect 306834 305368 306840 305380
rect 306432 305340 306840 305368
rect 306432 305328 306438 305340
rect 306834 305328 306840 305340
rect 306892 305328 306898 305380
rect 308030 305328 308036 305380
rect 308088 305368 308094 305380
rect 308766 305368 308772 305380
rect 308088 305340 308772 305368
rect 308088 305328 308094 305340
rect 308766 305328 308772 305340
rect 308824 305328 308830 305380
rect 309318 305328 309324 305380
rect 309376 305368 309382 305380
rect 309686 305368 309692 305380
rect 309376 305340 309692 305368
rect 309376 305328 309382 305340
rect 309686 305328 309692 305340
rect 309744 305328 309750 305380
rect 310514 305328 310520 305380
rect 310572 305368 310578 305380
rect 310882 305368 310888 305380
rect 310572 305340 310888 305368
rect 310572 305328 310578 305340
rect 310882 305328 310888 305340
rect 310940 305328 310946 305380
rect 311986 305328 311992 305380
rect 312044 305368 312050 305380
rect 313090 305368 313096 305380
rect 312044 305340 313096 305368
rect 312044 305328 312050 305340
rect 313090 305328 313096 305340
rect 313148 305328 313154 305380
rect 313550 305328 313556 305380
rect 313608 305368 313614 305380
rect 313826 305368 313832 305380
rect 313608 305340 313832 305368
rect 313608 305328 313614 305340
rect 313826 305328 313832 305340
rect 313884 305328 313890 305380
rect 314930 305328 314936 305380
rect 314988 305368 314994 305380
rect 315574 305368 315580 305380
rect 314988 305340 315580 305368
rect 314988 305328 314994 305340
rect 315574 305328 315580 305340
rect 315632 305328 315638 305380
rect 317690 305328 317696 305380
rect 317748 305368 317754 305380
rect 318518 305368 318524 305380
rect 317748 305340 318524 305368
rect 317748 305328 317754 305340
rect 318518 305328 318524 305340
rect 318576 305328 318582 305380
rect 318794 305328 318800 305380
rect 318852 305368 318858 305380
rect 319162 305368 319168 305380
rect 318852 305340 319168 305368
rect 318852 305328 318858 305340
rect 319162 305328 319168 305340
rect 319220 305328 319226 305380
rect 321554 305328 321560 305380
rect 321612 305368 321618 305380
rect 321922 305368 321928 305380
rect 321612 305340 321928 305368
rect 321612 305328 321618 305340
rect 321922 305328 321928 305340
rect 321980 305328 321986 305380
rect 323210 305328 323216 305380
rect 323268 305368 323274 305380
rect 323762 305368 323768 305380
rect 323268 305340 323768 305368
rect 323268 305328 323274 305340
rect 323762 305328 323768 305340
rect 323820 305328 323826 305380
rect 324406 305328 324412 305380
rect 324464 305368 324470 305380
rect 325142 305368 325148 305380
rect 324464 305340 325148 305368
rect 324464 305328 324470 305340
rect 325142 305328 325148 305340
rect 325200 305328 325206 305380
rect 325970 305328 325976 305380
rect 326028 305368 326034 305380
rect 326338 305368 326344 305380
rect 326028 305340 326344 305368
rect 326028 305328 326034 305340
rect 326338 305328 326344 305340
rect 326396 305328 326402 305380
rect 328638 305328 328644 305380
rect 328696 305368 328702 305380
rect 329006 305368 329012 305380
rect 328696 305340 329012 305368
rect 328696 305328 328702 305340
rect 329006 305328 329012 305340
rect 329064 305328 329070 305380
rect 330202 305328 330208 305380
rect 330260 305368 330266 305380
rect 331122 305368 331128 305380
rect 330260 305340 331128 305368
rect 330260 305328 330266 305340
rect 331122 305328 331128 305340
rect 331180 305328 331186 305380
rect 305086 305260 305092 305312
rect 305144 305300 305150 305312
rect 305914 305300 305920 305312
rect 305144 305272 305920 305300
rect 305144 305260 305150 305272
rect 305914 305260 305920 305272
rect 305972 305260 305978 305312
rect 308122 305260 308128 305312
rect 308180 305300 308186 305312
rect 308950 305300 308956 305312
rect 308180 305272 308956 305300
rect 308180 305260 308186 305272
rect 308950 305260 308956 305272
rect 309008 305260 309014 305312
rect 309226 305260 309232 305312
rect 309284 305300 309290 305312
rect 309502 305300 309508 305312
rect 309284 305272 309508 305300
rect 309284 305260 309290 305272
rect 309502 305260 309508 305272
rect 309560 305260 309566 305312
rect 314746 305260 314752 305312
rect 314804 305300 314810 305312
rect 315482 305300 315488 305312
rect 314804 305272 315488 305300
rect 314804 305260 314810 305272
rect 315482 305260 315488 305272
rect 315540 305260 315546 305312
rect 323026 305260 323032 305312
rect 323084 305300 323090 305312
rect 323946 305300 323952 305312
rect 323084 305272 323952 305300
rect 323084 305260 323090 305272
rect 323946 305260 323952 305272
rect 324004 305260 324010 305312
rect 326062 305260 326068 305312
rect 326120 305300 326126 305312
rect 326982 305300 326988 305312
rect 326120 305272 326988 305300
rect 326120 305260 326126 305272
rect 326982 305260 326988 305272
rect 327040 305260 327046 305312
rect 328730 305260 328736 305312
rect 328788 305300 328794 305312
rect 329374 305300 329380 305312
rect 328788 305272 329380 305300
rect 328788 305260 328794 305272
rect 329374 305260 329380 305272
rect 329432 305260 329438 305312
rect 330110 305260 330116 305312
rect 330168 305300 330174 305312
rect 330938 305300 330944 305312
rect 330168 305272 330944 305300
rect 330168 305260 330174 305272
rect 330938 305260 330944 305272
rect 330996 305260 331002 305312
rect 298060 305204 302234 305232
rect 298060 305192 298066 305204
rect 306374 305192 306380 305244
rect 306432 305232 306438 305244
rect 307294 305232 307300 305244
rect 306432 305204 307300 305232
rect 306432 305192 306438 305204
rect 307294 305192 307300 305204
rect 307352 305192 307358 305244
rect 310514 305192 310520 305244
rect 310572 305232 310578 305244
rect 311342 305232 311348 305244
rect 310572 305204 311348 305232
rect 310572 305192 310578 305204
rect 311342 305192 311348 305204
rect 311400 305192 311406 305244
rect 314654 305192 314660 305244
rect 314712 305232 314718 305244
rect 315942 305232 315948 305244
rect 314712 305204 315948 305232
rect 314712 305192 314718 305204
rect 315942 305192 315948 305204
rect 316000 305192 316006 305244
rect 321554 305192 321560 305244
rect 321612 305232 321618 305244
rect 322658 305232 322664 305244
rect 321612 305204 322664 305232
rect 321612 305192 321618 305204
rect 322658 305192 322664 305204
rect 322716 305192 322722 305244
rect 328546 305192 328552 305244
rect 328604 305232 328610 305244
rect 329466 305232 329472 305244
rect 328604 305204 329472 305232
rect 328604 305192 328610 305204
rect 329466 305192 329472 305204
rect 329524 305192 329530 305244
rect 329926 305192 329932 305244
rect 329984 305232 329990 305244
rect 330570 305232 330576 305244
rect 329984 305204 330576 305232
rect 329984 305192 329990 305204
rect 330570 305192 330576 305204
rect 330628 305192 330634 305244
rect 331232 305164 331260 305408
rect 332502 305396 332508 305448
rect 332560 305436 332566 305448
rect 338758 305436 338764 305448
rect 332560 305408 338764 305436
rect 332560 305396 332566 305408
rect 338758 305396 338764 305408
rect 338816 305396 338822 305448
rect 343634 305436 343640 305448
rect 340846 305408 343640 305436
rect 331398 305328 331404 305380
rect 331456 305368 331462 305380
rect 332226 305368 332232 305380
rect 331456 305340 332232 305368
rect 331456 305328 331462 305340
rect 332226 305328 332232 305340
rect 332284 305328 332290 305380
rect 332778 305328 332784 305380
rect 332836 305368 332842 305380
rect 333514 305368 333520 305380
rect 332836 305340 333520 305368
rect 332836 305328 332842 305340
rect 333514 305328 333520 305340
rect 333572 305328 333578 305380
rect 331950 305260 331956 305312
rect 332008 305300 332014 305312
rect 339862 305300 339868 305312
rect 332008 305272 339868 305300
rect 332008 305260 332014 305272
rect 339862 305260 339868 305272
rect 339920 305260 339926 305312
rect 340846 305164 340874 305408
rect 343634 305396 343640 305408
rect 343692 305396 343698 305448
rect 331232 305136 340874 305164
rect 254026 304784 254032 304836
rect 254084 304824 254090 304836
rect 254302 304824 254308 304836
rect 254084 304796 254308 304824
rect 254084 304784 254090 304796
rect 254302 304784 254308 304796
rect 254360 304784 254366 304836
rect 254026 304648 254032 304700
rect 254084 304688 254090 304700
rect 254486 304688 254492 304700
rect 254084 304660 254492 304688
rect 254084 304648 254090 304660
rect 254486 304648 254492 304660
rect 254544 304648 254550 304700
rect 316586 304444 316592 304496
rect 316644 304484 316650 304496
rect 443638 304484 443644 304496
rect 316644 304456 443644 304484
rect 316644 304444 316650 304456
rect 443638 304444 443644 304456
rect 443696 304444 443702 304496
rect 85574 304376 85580 304428
rect 85632 304416 85638 304428
rect 245654 304416 245660 304428
rect 85632 304388 245660 304416
rect 85632 304376 85638 304388
rect 245654 304376 245660 304388
rect 245712 304376 245718 304428
rect 319622 304376 319628 304428
rect 319680 304416 319686 304428
rect 485038 304416 485044 304428
rect 319680 304388 485044 304416
rect 319680 304376 319686 304388
rect 485038 304376 485044 304388
rect 485096 304376 485102 304428
rect 82170 304308 82176 304360
rect 82228 304348 82234 304360
rect 244366 304348 244372 304360
rect 82228 304320 244372 304348
rect 82228 304308 82234 304320
rect 244366 304308 244372 304320
rect 244424 304308 244430 304360
rect 325510 304308 325516 304360
rect 325568 304348 325574 304360
rect 516778 304348 516784 304360
rect 325568 304320 516784 304348
rect 325568 304308 325574 304320
rect 516778 304308 516784 304320
rect 516836 304308 516842 304360
rect 7558 304240 7564 304292
rect 7616 304280 7622 304292
rect 230474 304280 230480 304292
rect 7616 304252 230480 304280
rect 7616 304240 7622 304252
rect 230474 304240 230480 304252
rect 230532 304240 230538 304292
rect 233418 304240 233424 304292
rect 233476 304280 233482 304292
rect 233602 304280 233608 304292
rect 233476 304252 233608 304280
rect 233476 304240 233482 304252
rect 233602 304240 233608 304252
rect 233660 304240 233666 304292
rect 256970 304240 256976 304292
rect 257028 304280 257034 304292
rect 257246 304280 257252 304292
rect 257028 304252 257252 304280
rect 257028 304240 257034 304252
rect 257246 304240 257252 304252
rect 257304 304240 257310 304292
rect 276290 304240 276296 304292
rect 276348 304280 276354 304292
rect 276566 304280 276572 304292
rect 276348 304252 276572 304280
rect 276348 304240 276354 304252
rect 276566 304240 276572 304252
rect 276624 304240 276630 304292
rect 304902 304240 304908 304292
rect 304960 304280 304966 304292
rect 305454 304280 305460 304292
rect 304960 304252 305460 304280
rect 304960 304240 304966 304252
rect 305454 304240 305460 304252
rect 305512 304240 305518 304292
rect 310790 304240 310796 304292
rect 310848 304280 310854 304292
rect 311158 304280 311164 304292
rect 310848 304252 311164 304280
rect 310848 304240 310854 304252
rect 311158 304240 311164 304252
rect 311216 304240 311222 304292
rect 313642 304240 313648 304292
rect 313700 304280 313706 304292
rect 313918 304280 313924 304292
rect 313700 304252 313924 304280
rect 313700 304240 313706 304252
rect 313918 304240 313924 304252
rect 313976 304240 313982 304292
rect 318978 304240 318984 304292
rect 319036 304280 319042 304292
rect 319254 304280 319260 304292
rect 319036 304252 319260 304280
rect 319036 304240 319042 304252
rect 319254 304240 319260 304252
rect 319312 304240 319318 304292
rect 334526 304240 334532 304292
rect 334584 304280 334590 304292
rect 563698 304280 563704 304292
rect 334584 304252 563704 304280
rect 334584 304240 334590 304252
rect 563698 304240 563704 304252
rect 563756 304240 563762 304292
rect 291378 304172 291384 304224
rect 291436 304212 291442 304224
rect 292298 304212 292304 304224
rect 291436 304184 292304 304212
rect 291436 304172 291442 304184
rect 292298 304172 292304 304184
rect 292356 304172 292362 304224
rect 230658 304104 230664 304156
rect 230716 304144 230722 304156
rect 231762 304144 231768 304156
rect 230716 304116 231768 304144
rect 230716 304104 230722 304116
rect 231762 304104 231768 304116
rect 231820 304104 231826 304156
rect 248598 304104 248604 304156
rect 248656 304144 248662 304156
rect 249610 304144 249616 304156
rect 248656 304116 249616 304144
rect 248656 304104 248662 304116
rect 249610 304104 249616 304116
rect 249668 304104 249674 304156
rect 251542 303968 251548 304020
rect 251600 304008 251606 304020
rect 252462 304008 252468 304020
rect 251600 303980 252468 304008
rect 251600 303968 251606 303980
rect 252462 303968 252468 303980
rect 252520 303968 252526 304020
rect 273438 303968 273444 304020
rect 273496 304008 273502 304020
rect 274266 304008 274272 304020
rect 273496 303980 274272 304008
rect 273496 303968 273502 303980
rect 274266 303968 274272 303980
rect 274324 303968 274330 304020
rect 318794 303696 318800 303748
rect 318852 303736 318858 303748
rect 319898 303736 319904 303748
rect 318852 303708 319904 303736
rect 318852 303696 318858 303708
rect 319898 303696 319904 303708
rect 319956 303696 319962 303748
rect 275922 303560 275928 303612
rect 275980 303600 275986 303612
rect 341242 303600 341248 303612
rect 275980 303572 341248 303600
rect 275980 303560 275986 303572
rect 341242 303560 341248 303572
rect 341300 303560 341306 303612
rect 272518 303492 272524 303544
rect 272576 303532 272582 303544
rect 342346 303532 342352 303544
rect 272576 303504 342352 303532
rect 272576 303492 272582 303504
rect 342346 303492 342352 303504
rect 342404 303492 342410 303544
rect 264974 303424 264980 303476
rect 265032 303464 265038 303476
rect 265894 303464 265900 303476
rect 265032 303436 265900 303464
rect 265032 303424 265038 303436
rect 265894 303424 265900 303436
rect 265952 303424 265958 303476
rect 272794 303424 272800 303476
rect 272852 303464 272858 303476
rect 343726 303464 343732 303476
rect 272852 303436 343732 303464
rect 272852 303424 272858 303436
rect 343726 303424 343732 303436
rect 343784 303424 343790 303476
rect 269850 303356 269856 303408
rect 269908 303396 269914 303408
rect 344830 303396 344836 303408
rect 269908 303368 344836 303396
rect 269908 303356 269914 303368
rect 344830 303356 344836 303368
rect 344888 303356 344894 303408
rect 279878 303288 279884 303340
rect 279936 303328 279942 303340
rect 355134 303328 355140 303340
rect 279936 303300 355140 303328
rect 279936 303288 279942 303300
rect 355134 303288 355140 303300
rect 355192 303288 355198 303340
rect 269942 303220 269948 303272
rect 270000 303260 270006 303272
rect 345106 303260 345112 303272
rect 270000 303232 345112 303260
rect 270000 303220 270006 303232
rect 345106 303220 345112 303232
rect 345164 303220 345170 303272
rect 270034 303152 270040 303204
rect 270092 303192 270098 303204
rect 346394 303192 346400 303204
rect 270092 303164 346400 303192
rect 270092 303152 270098 303164
rect 346394 303152 346400 303164
rect 346452 303152 346458 303204
rect 278130 303084 278136 303136
rect 278188 303124 278194 303136
rect 357526 303124 357532 303136
rect 278188 303096 357532 303124
rect 278188 303084 278194 303096
rect 357526 303084 357532 303096
rect 357584 303084 357590 303136
rect 93118 303016 93124 303068
rect 93176 303056 93182 303068
rect 245102 303056 245108 303068
rect 93176 303028 245108 303056
rect 93176 303016 93182 303028
rect 245102 303016 245108 303028
rect 245160 303016 245166 303068
rect 276106 303016 276112 303068
rect 276164 303056 276170 303068
rect 277210 303056 277216 303068
rect 276164 303028 277216 303056
rect 276164 303016 276170 303028
rect 277210 303016 277216 303028
rect 277268 303016 277274 303068
rect 278222 303016 278228 303068
rect 278280 303056 278286 303068
rect 358906 303056 358912 303068
rect 278280 303028 358912 303056
rect 278280 303016 278286 303028
rect 358906 303016 358912 303028
rect 358964 303016 358970 303068
rect 93854 302948 93860 303000
rect 93912 302988 93918 303000
rect 247218 302988 247224 303000
rect 93912 302960 247224 302988
rect 93912 302948 93918 302960
rect 247218 302948 247224 302960
rect 247276 302948 247282 303000
rect 275370 302948 275376 303000
rect 275428 302988 275434 303000
rect 358814 302988 358820 303000
rect 275428 302960 358820 302988
rect 275428 302948 275434 302960
rect 358814 302948 358820 302960
rect 358872 302948 358878 303000
rect 8938 302880 8944 302932
rect 8996 302920 9002 302932
rect 231394 302920 231400 302932
rect 8996 302892 231400 302920
rect 8996 302880 9002 302892
rect 231394 302880 231400 302892
rect 231452 302880 231458 302932
rect 275462 302880 275468 302932
rect 275520 302920 275526 302932
rect 359090 302920 359096 302932
rect 275520 302892 359096 302920
rect 275520 302880 275526 302892
rect 359090 302880 359096 302892
rect 359148 302880 359154 302932
rect 277118 302812 277124 302864
rect 277176 302852 277182 302864
rect 277302 302852 277308 302864
rect 277176 302824 277308 302852
rect 277176 302812 277182 302824
rect 277302 302812 277308 302824
rect 277360 302812 277366 302864
rect 293770 302812 293776 302864
rect 293828 302852 293834 302864
rect 342806 302852 342812 302864
rect 293828 302824 342812 302852
rect 293828 302812 293834 302824
rect 342806 302812 342812 302824
rect 342864 302812 342870 302864
rect 263594 302744 263600 302796
rect 263652 302784 263658 302796
rect 264606 302784 264612 302796
rect 263652 302756 264612 302784
rect 263652 302744 263658 302756
rect 264606 302744 264612 302756
rect 264664 302744 264670 302796
rect 294966 302744 294972 302796
rect 295024 302784 295030 302796
rect 342530 302784 342536 302796
rect 295024 302756 342536 302784
rect 295024 302744 295030 302756
rect 342530 302744 342536 302756
rect 342588 302744 342594 302796
rect 293586 302676 293592 302728
rect 293644 302716 293650 302728
rect 338114 302716 338120 302728
rect 293644 302688 338120 302716
rect 293644 302676 293650 302688
rect 338114 302676 338120 302688
rect 338172 302676 338178 302728
rect 258258 302608 258264 302660
rect 258316 302648 258322 302660
rect 258534 302648 258540 302660
rect 258316 302620 258540 302648
rect 258316 302608 258322 302620
rect 258534 302608 258540 302620
rect 258592 302608 258598 302660
rect 320542 301588 320548 301640
rect 320600 301628 320606 301640
rect 491938 301628 491944 301640
rect 320600 301600 491944 301628
rect 320600 301588 320606 301600
rect 491938 301588 491944 301600
rect 491996 301588 492002 301640
rect 48958 301520 48964 301572
rect 49016 301560 49022 301572
rect 239122 301560 239128 301572
rect 49016 301532 239128 301560
rect 49016 301520 49022 301532
rect 239122 301520 239128 301532
rect 239180 301520 239186 301572
rect 328914 301520 328920 301572
rect 328972 301560 328978 301572
rect 534718 301560 534724 301572
rect 328972 301532 534724 301560
rect 328972 301520 328978 301532
rect 534718 301520 534724 301532
rect 534776 301520 534782 301572
rect 43438 301452 43444 301504
rect 43496 301492 43502 301504
rect 237374 301492 237380 301504
rect 43496 301464 237380 301492
rect 43496 301452 43502 301464
rect 237374 301452 237380 301464
rect 237432 301452 237438 301504
rect 334802 301452 334808 301504
rect 334860 301492 334866 301504
rect 565814 301492 565820 301504
rect 334860 301464 565820 301492
rect 334860 301452 334866 301464
rect 565814 301452 565820 301464
rect 565872 301452 565878 301504
rect 285214 300772 285220 300824
rect 285272 300812 285278 300824
rect 336918 300812 336924 300824
rect 285272 300784 336924 300812
rect 285272 300772 285278 300784
rect 336918 300772 336924 300784
rect 336976 300772 336982 300824
rect 285398 300704 285404 300756
rect 285456 300744 285462 300756
rect 338298 300744 338304 300756
rect 285456 300716 338304 300744
rect 285456 300704 285462 300716
rect 338298 300704 338304 300716
rect 338356 300704 338362 300756
rect 290826 300636 290832 300688
rect 290884 300676 290890 300688
rect 345014 300676 345020 300688
rect 290884 300648 345020 300676
rect 290884 300636 290890 300648
rect 345014 300636 345020 300648
rect 345072 300636 345078 300688
rect 286962 300568 286968 300620
rect 287020 300608 287026 300620
rect 346578 300608 346584 300620
rect 287020 300580 346584 300608
rect 287020 300568 287026 300580
rect 346578 300568 346584 300580
rect 346636 300568 346642 300620
rect 267918 300500 267924 300552
rect 267976 300540 267982 300552
rect 268286 300540 268292 300552
rect 267976 300512 268292 300540
rect 267976 300500 267982 300512
rect 268286 300500 268292 300512
rect 268344 300500 268350 300552
rect 296622 300500 296628 300552
rect 296680 300540 296686 300552
rect 357618 300540 357624 300552
rect 296680 300512 357624 300540
rect 296680 300500 296686 300512
rect 357618 300500 357624 300512
rect 357676 300500 357682 300552
rect 241882 300432 241888 300484
rect 241940 300472 241946 300484
rect 242066 300472 242072 300484
rect 241940 300444 242072 300472
rect 241940 300432 241946 300444
rect 242066 300432 242072 300444
rect 242124 300432 242130 300484
rect 283834 300432 283840 300484
rect 283892 300472 283898 300484
rect 345290 300472 345296 300484
rect 283892 300444 345296 300472
rect 283892 300432 283898 300444
rect 345290 300432 345296 300444
rect 345348 300432 345354 300484
rect 282546 300364 282552 300416
rect 282604 300404 282610 300416
rect 347314 300404 347320 300416
rect 282604 300376 347320 300404
rect 282604 300364 282610 300376
rect 347314 300364 347320 300376
rect 347372 300364 347378 300416
rect 285490 300296 285496 300348
rect 285548 300336 285554 300348
rect 351086 300336 351092 300348
rect 285548 300308 351092 300336
rect 285548 300296 285554 300308
rect 351086 300296 351092 300308
rect 351144 300296 351150 300348
rect 292298 300228 292304 300280
rect 292356 300268 292362 300280
rect 357894 300268 357900 300280
rect 292356 300240 357900 300268
rect 292356 300228 292362 300240
rect 357894 300228 357900 300240
rect 357952 300228 357958 300280
rect 53098 300160 53104 300212
rect 53156 300200 53162 300212
rect 238846 300200 238852 300212
rect 53156 300172 238852 300200
rect 53156 300160 53162 300172
rect 238846 300160 238852 300172
rect 238904 300160 238910 300212
rect 279602 300160 279608 300212
rect 279660 300200 279666 300212
rect 349338 300200 349344 300212
rect 279660 300172 349344 300200
rect 279660 300160 279666 300172
rect 349338 300160 349344 300172
rect 349396 300160 349402 300212
rect 10318 300092 10324 300144
rect 10376 300132 10382 300144
rect 231026 300132 231032 300144
rect 10376 300104 231032 300132
rect 10376 300092 10382 300104
rect 231026 300092 231032 300104
rect 231084 300092 231090 300144
rect 285306 300092 285312 300144
rect 285364 300132 285370 300144
rect 360194 300132 360200 300144
rect 285364 300104 360200 300132
rect 285364 300092 285370 300104
rect 360194 300092 360200 300104
rect 360252 300092 360258 300144
rect 286870 300024 286876 300076
rect 286928 300064 286934 300076
rect 338206 300064 338212 300076
rect 286928 300036 338212 300064
rect 286928 300024 286934 300036
rect 338206 300024 338212 300036
rect 338264 300024 338270 300076
rect 288250 299956 288256 300008
rect 288308 299996 288314 300008
rect 340506 299996 340512 300008
rect 288308 299968 340512 299996
rect 288308 299956 288314 299968
rect 340506 299956 340512 299968
rect 340564 299956 340570 300008
rect 290734 299888 290740 299940
rect 290792 299928 290798 299940
rect 341426 299928 341432 299940
rect 290792 299900 341432 299928
rect 290792 299888 290798 299900
rect 341426 299888 341432 299900
rect 341484 299888 341490 299940
rect 313734 298936 313740 298988
rect 313792 298976 313798 298988
rect 454034 298976 454040 298988
rect 313792 298948 454040 298976
rect 313792 298936 313798 298948
rect 454034 298936 454040 298948
rect 454092 298936 454098 298988
rect 323394 298868 323400 298920
rect 323452 298908 323458 298920
rect 502978 298908 502984 298920
rect 323452 298880 502984 298908
rect 323452 298868 323458 298880
rect 502978 298868 502984 298880
rect 503036 298868 503042 298920
rect 326246 298800 326252 298852
rect 326304 298840 326310 298852
rect 520274 298840 520280 298852
rect 326304 298812 520280 298840
rect 326304 298800 326310 298812
rect 520274 298800 520280 298812
rect 520332 298800 520338 298852
rect 53834 298732 53840 298784
rect 53892 298772 53898 298784
rect 238754 298772 238760 298784
rect 53892 298744 238760 298772
rect 53892 298732 53898 298744
rect 238754 298732 238760 298744
rect 238812 298732 238818 298784
rect 333054 298732 333060 298784
rect 333112 298772 333118 298784
rect 557534 298772 557540 298784
rect 333112 298744 557540 298772
rect 333112 298732 333118 298744
rect 557534 298732 557540 298744
rect 557592 298732 557598 298784
rect 251174 298596 251180 298648
rect 251232 298636 251238 298648
rect 251358 298636 251364 298648
rect 251232 298608 251364 298636
rect 251232 298596 251238 298608
rect 251358 298596 251364 298608
rect 251416 298596 251422 298648
rect 278590 297780 278596 297832
rect 278648 297820 278654 297832
rect 338390 297820 338396 297832
rect 278648 297792 338396 297820
rect 278648 297780 278654 297792
rect 338390 297780 338396 297792
rect 338448 297780 338454 297832
rect 282454 297712 282460 297764
rect 282512 297752 282518 297764
rect 343818 297752 343824 297764
rect 282512 297724 343824 297752
rect 282512 297712 282518 297724
rect 343818 297712 343824 297724
rect 343876 297712 343882 297764
rect 275830 297644 275836 297696
rect 275888 297684 275894 297696
rect 339678 297684 339684 297696
rect 275888 297656 339684 297684
rect 275888 297644 275894 297656
rect 339678 297644 339684 297656
rect 339736 297644 339742 297696
rect 283926 297576 283932 297628
rect 283984 297616 283990 297628
rect 358998 297616 359004 297628
rect 283984 297588 359004 297616
rect 283984 297576 283990 297588
rect 358998 297576 359004 297588
rect 359056 297576 359062 297628
rect 323302 297508 323308 297560
rect 323360 297548 323366 297560
rect 507854 297548 507860 297560
rect 323360 297520 507860 297548
rect 323360 297508 323366 297520
rect 507854 297508 507860 297520
rect 507912 297508 507918 297560
rect 86954 297440 86960 297492
rect 87012 297480 87018 297492
rect 245930 297480 245936 297492
rect 87012 297452 245936 297480
rect 87012 297440 87018 297452
rect 245930 297440 245936 297452
rect 245988 297440 245994 297492
rect 269574 297440 269580 297492
rect 269632 297440 269638 297492
rect 285858 297440 285864 297492
rect 285916 297440 285922 297492
rect 332962 297440 332968 297492
rect 333020 297480 333026 297492
rect 560294 297480 560300 297492
rect 333020 297452 560300 297480
rect 333020 297440 333026 297452
rect 560294 297440 560300 297452
rect 560352 297440 560358 297492
rect 60734 297372 60740 297424
rect 60792 297412 60798 297424
rect 240410 297412 240416 297424
rect 60792 297384 240416 297412
rect 60792 297372 60798 297384
rect 240410 297372 240416 297384
rect 240468 297372 240474 297424
rect 269592 297288 269620 297440
rect 269574 297236 269580 297288
rect 269632 297236 269638 297288
rect 285876 297276 285904 297440
rect 334250 297372 334256 297424
rect 334308 297412 334314 297424
rect 570598 297412 570604 297424
rect 334308 297384 570604 297412
rect 334308 297372 334314 297384
rect 570598 297372 570604 297384
rect 570656 297372 570662 297424
rect 285950 297276 285956 297288
rect 285876 297248 285956 297276
rect 285950 297236 285956 297248
rect 286008 297236 286014 297288
rect 93946 296012 93952 296064
rect 94004 296052 94010 296064
rect 247586 296052 247592 296064
rect 94004 296024 247592 296052
rect 94004 296012 94010 296024
rect 247586 296012 247592 296024
rect 247644 296012 247650 296064
rect 316310 296012 316316 296064
rect 316368 296052 316374 296064
rect 467098 296052 467104 296064
rect 316368 296024 467104 296052
rect 316368 296012 316374 296024
rect 467098 296012 467104 296024
rect 467156 296012 467162 296064
rect 66898 295944 66904 295996
rect 66956 295984 66962 295996
rect 241974 295984 241980 295996
rect 66956 295956 241980 295984
rect 66956 295944 66962 295956
rect 241974 295944 241980 295956
rect 242032 295944 242038 295996
rect 324682 295944 324688 295996
rect 324740 295984 324746 295996
rect 514018 295984 514024 295996
rect 324740 295956 514024 295984
rect 324740 295944 324746 295956
rect 514018 295944 514024 295956
rect 514076 295944 514082 295996
rect 316218 294720 316224 294772
rect 316276 294760 316282 294772
rect 471238 294760 471244 294772
rect 316276 294732 471244 294760
rect 316276 294720 316282 294732
rect 471238 294720 471244 294732
rect 471296 294720 471302 294772
rect 69014 294652 69020 294704
rect 69072 294692 69078 294704
rect 241790 294692 241796 294704
rect 69072 294664 241796 294692
rect 69072 294652 69078 294664
rect 241790 294652 241796 294664
rect 241848 294652 241854 294704
rect 327534 294652 327540 294704
rect 327592 294692 327598 294704
rect 529934 294692 529940 294704
rect 327592 294664 529940 294692
rect 327592 294652 327598 294664
rect 529934 294652 529940 294664
rect 529992 294652 529998 294704
rect 31018 294584 31024 294636
rect 31076 294624 31082 294636
rect 234890 294624 234896 294636
rect 31076 294596 234896 294624
rect 31076 294584 31082 294596
rect 234890 294584 234896 294596
rect 234948 294584 234954 294636
rect 283098 294584 283104 294636
rect 283156 294624 283162 294636
rect 283282 294624 283288 294636
rect 283156 294596 283288 294624
rect 283156 294584 283162 294596
rect 283282 294584 283288 294596
rect 283340 294584 283346 294636
rect 328822 294584 328828 294636
rect 328880 294624 328886 294636
rect 535454 294624 535460 294636
rect 328880 294596 535460 294624
rect 328880 294584 328886 294596
rect 535454 294584 535460 294596
rect 535512 294584 535518 294636
rect 3326 293904 3332 293956
rect 3384 293944 3390 293956
rect 228450 293944 228456 293956
rect 3384 293916 228456 293944
rect 3384 293904 3390 293916
rect 228450 293904 228456 293916
rect 228508 293904 228514 293956
rect 54478 293224 54484 293276
rect 54536 293264 54542 293276
rect 239030 293264 239036 293276
rect 54536 293236 239036 293264
rect 54536 293224 54542 293236
rect 239030 293224 239036 293236
rect 239088 293224 239094 293276
rect 327442 293224 327448 293276
rect 327500 293264 327506 293276
rect 527818 293264 527824 293276
rect 327500 293236 527824 293264
rect 327500 293224 327506 293236
rect 527818 293224 527824 293236
rect 527876 293224 527882 293276
rect 71774 291864 71780 291916
rect 71832 291904 71838 291916
rect 243078 291904 243084 291916
rect 71832 291876 243084 291904
rect 71832 291864 71838 291876
rect 243078 291864 243084 291876
rect 243136 291864 243142 291916
rect 34514 291796 34520 291848
rect 34572 291836 34578 291848
rect 236270 291836 236276 291848
rect 34572 291808 236276 291836
rect 34572 291796 34578 291808
rect 236270 291796 236276 291808
rect 236328 291796 236334 291848
rect 328730 291796 328736 291848
rect 328788 291836 328794 291848
rect 538858 291836 538864 291848
rect 328788 291808 538864 291836
rect 328788 291796 328794 291808
rect 538858 291796 538864 291808
rect 538916 291796 538922 291848
rect 269482 291116 269488 291168
rect 269540 291156 269546 291168
rect 269666 291156 269672 291168
rect 269540 291128 269672 291156
rect 269540 291116 269546 291128
rect 269666 291116 269672 291128
rect 269724 291116 269730 291168
rect 331674 290504 331680 290556
rect 331732 290544 331738 290556
rect 549898 290544 549904 290556
rect 331732 290516 549904 290544
rect 331732 290504 331738 290516
rect 549898 290504 549904 290516
rect 549956 290504 549962 290556
rect 41414 290436 41420 290488
rect 41472 290476 41478 290488
rect 237650 290476 237656 290488
rect 41472 290448 237656 290476
rect 41472 290436 41478 290448
rect 237650 290436 237656 290448
rect 237708 290436 237714 290488
rect 334158 290436 334164 290488
rect 334216 290476 334222 290488
rect 567194 290476 567200 290488
rect 334216 290448 567200 290476
rect 334216 290436 334222 290448
rect 567194 290436 567200 290448
rect 567252 290436 567258 290488
rect 58618 289144 58624 289196
rect 58676 289184 58682 289196
rect 240318 289184 240324 289196
rect 58676 289156 240324 289184
rect 58676 289144 58682 289156
rect 240318 289144 240324 289156
rect 240376 289144 240382 289196
rect 331582 289144 331588 289196
rect 331640 289184 331646 289196
rect 552658 289184 552664 289196
rect 331640 289156 552664 289184
rect 331640 289144 331646 289156
rect 552658 289144 552664 289156
rect 552716 289144 552722 289196
rect 13078 289076 13084 289128
rect 13136 289116 13142 289128
rect 232130 289116 232136 289128
rect 13136 289088 232136 289116
rect 13136 289076 13142 289088
rect 232130 289076 232136 289088
rect 232188 289076 232194 289128
rect 334066 289076 334072 289128
rect 334124 289116 334130 289128
rect 567838 289116 567844 289128
rect 334124 289088 567844 289116
rect 334124 289076 334130 289088
rect 567838 289076 567844 289088
rect 567896 289076 567902 289128
rect 312170 287784 312176 287836
rect 312228 287824 312234 287836
rect 448514 287824 448520 287836
rect 312228 287796 448520 287824
rect 312228 287784 312234 287796
rect 448514 287784 448520 287796
rect 448572 287784 448578 287836
rect 312262 287716 312268 287768
rect 312320 287756 312326 287768
rect 449894 287756 449900 287768
rect 312320 287728 449900 287756
rect 312320 287716 312326 287728
rect 449894 287716 449900 287728
rect 449952 287716 449958 287768
rect 9674 287648 9680 287700
rect 9732 287688 9738 287700
rect 230658 287688 230664 287700
rect 9732 287660 230664 287688
rect 9732 287648 9738 287660
rect 230658 287648 230664 287660
rect 230716 287648 230722 287700
rect 332870 287648 332876 287700
rect 332928 287688 332934 287700
rect 561674 287688 561680 287700
rect 332928 287660 561680 287688
rect 332928 287648 332934 287660
rect 561674 287648 561680 287660
rect 561732 287648 561738 287700
rect 315114 286492 315120 286544
rect 315172 286532 315178 286544
rect 462314 286532 462320 286544
rect 315172 286504 462320 286532
rect 315172 286492 315178 286504
rect 462314 286492 462320 286504
rect 462372 286492 462378 286544
rect 318150 286424 318156 286476
rect 318208 286464 318214 286476
rect 467834 286464 467840 286476
rect 318208 286436 467840 286464
rect 318208 286424 318214 286436
rect 467834 286424 467840 286436
rect 467892 286424 467898 286476
rect 89714 286356 89720 286408
rect 89772 286396 89778 286408
rect 245838 286396 245844 286408
rect 89772 286368 245844 286396
rect 89772 286356 89778 286368
rect 245838 286356 245844 286368
rect 245896 286356 245902 286408
rect 319162 286356 319168 286408
rect 319220 286396 319226 286408
rect 481634 286396 481640 286408
rect 319220 286368 481640 286396
rect 319220 286356 319226 286368
rect 481634 286356 481640 286368
rect 481692 286356 481698 286408
rect 46290 286288 46296 286340
rect 46348 286328 46354 286340
rect 237558 286328 237564 286340
rect 46348 286300 237564 286328
rect 46348 286288 46354 286300
rect 237558 286288 237564 286300
rect 237616 286288 237622 286340
rect 335814 286288 335820 286340
rect 335872 286328 335878 286340
rect 575474 286328 575480 286340
rect 335872 286300 575480 286328
rect 335872 286288 335878 286300
rect 575474 286288 575480 286300
rect 575532 286288 575538 286340
rect 96614 284996 96620 285048
rect 96672 285036 96678 285048
rect 247310 285036 247316 285048
rect 96672 285008 247316 285036
rect 96672 284996 96678 285008
rect 247310 284996 247316 285008
rect 247368 284996 247374 285048
rect 39390 284928 39396 284980
rect 39448 284968 39454 284980
rect 236178 284968 236184 284980
rect 39448 284940 236184 284968
rect 39448 284928 39454 284940
rect 236178 284928 236184 284940
rect 236236 284928 236242 284980
rect 313642 284928 313648 284980
rect 313700 284968 313706 284980
rect 453298 284968 453304 284980
rect 313700 284940 453304 284968
rect 313700 284928 313706 284940
rect 453298 284928 453304 284940
rect 453356 284928 453362 284980
rect 313550 283704 313556 283756
rect 313608 283744 313614 283756
rect 456794 283744 456800 283756
rect 313608 283716 456800 283744
rect 313608 283704 313614 283716
rect 456794 283704 456800 283716
rect 456852 283704 456858 283756
rect 67634 283636 67640 283688
rect 67692 283676 67698 283688
rect 241698 283676 241704 283688
rect 67692 283648 241704 283676
rect 67692 283636 67698 283648
rect 241698 283636 241704 283648
rect 241756 283636 241762 283688
rect 317690 283636 317696 283688
rect 317748 283676 317754 283688
rect 481726 283676 481732 283688
rect 317748 283648 481732 283676
rect 317748 283636 317754 283648
rect 481726 283636 481732 283648
rect 481784 283636 481790 283688
rect 16574 283568 16580 283620
rect 16632 283608 16638 283620
rect 232038 283608 232044 283620
rect 16632 283580 232044 283608
rect 16632 283568 16638 283580
rect 232038 283568 232044 283580
rect 232096 283568 232102 283620
rect 333974 283568 333980 283620
rect 334032 283608 334038 283620
rect 571334 283608 571340 283620
rect 334032 283580 571340 283608
rect 334032 283568 334038 283580
rect 571334 283568 571340 283580
rect 571392 283568 571398 283620
rect 318058 282276 318064 282328
rect 318116 282316 318122 282328
rect 460934 282316 460940 282328
rect 318116 282288 460940 282316
rect 318116 282276 318122 282288
rect 460934 282276 460940 282288
rect 460992 282276 460998 282328
rect 74534 282208 74540 282260
rect 74592 282248 74598 282260
rect 235258 282248 235264 282260
rect 74592 282220 235264 282248
rect 74592 282208 74598 282220
rect 235258 282208 235264 282220
rect 235316 282208 235322 282260
rect 315022 282208 315028 282260
rect 315080 282248 315086 282260
rect 459554 282248 459560 282260
rect 315080 282220 459560 282248
rect 315080 282208 315086 282220
rect 459554 282208 459560 282220
rect 459612 282208 459618 282260
rect 20714 282140 20720 282192
rect 20772 282180 20778 282192
rect 233602 282180 233608 282192
rect 20772 282152 233608 282180
rect 20772 282140 20778 282152
rect 233602 282140 233608 282152
rect 233660 282140 233666 282192
rect 319070 282140 319076 282192
rect 319128 282180 319134 282192
rect 484394 282180 484400 282192
rect 319128 282152 484400 282180
rect 319128 282140 319134 282152
rect 484394 282140 484400 282152
rect 484452 282140 484458 282192
rect 320818 280916 320824 280968
rect 320876 280956 320882 280968
rect 474734 280956 474740 280968
rect 320876 280928 474740 280956
rect 320876 280916 320882 280928
rect 474734 280916 474740 280928
rect 474792 280916 474798 280968
rect 88978 280848 88984 280900
rect 89036 280888 89042 280900
rect 245746 280888 245752 280900
rect 89036 280860 245752 280888
rect 89036 280848 89042 280860
rect 245746 280848 245752 280860
rect 245804 280848 245810 280900
rect 316126 280848 316132 280900
rect 316184 280888 316190 280900
rect 472618 280888 472624 280900
rect 316184 280860 472624 280888
rect 316184 280848 316190 280860
rect 472618 280848 472624 280860
rect 472676 280848 472682 280900
rect 26234 280780 26240 280832
rect 26292 280820 26298 280832
rect 234798 280820 234804 280832
rect 26292 280792 234804 280820
rect 26292 280780 26298 280792
rect 234798 280780 234804 280792
rect 234856 280780 234862 280832
rect 321830 280780 321836 280832
rect 321888 280820 321894 280832
rect 502334 280820 502340 280832
rect 321888 280792 502340 280820
rect 321888 280780 321894 280792
rect 502334 280780 502340 280792
rect 502392 280780 502398 280832
rect 92474 279488 92480 279540
rect 92532 279528 92538 279540
rect 247218 279528 247224 279540
rect 92532 279500 247224 279528
rect 92532 279488 92538 279500
rect 247218 279488 247224 279500
rect 247276 279488 247282 279540
rect 318978 279488 318984 279540
rect 319036 279528 319042 279540
rect 485774 279528 485780 279540
rect 319036 279500 485780 279528
rect 319036 279488 319042 279500
rect 485774 279488 485780 279500
rect 485832 279488 485838 279540
rect 40678 279420 40684 279472
rect 40736 279460 40742 279472
rect 234706 279460 234712 279472
rect 40736 279432 234712 279460
rect 40736 279420 40742 279432
rect 234706 279420 234712 279432
rect 234764 279420 234770 279472
rect 324590 279420 324596 279472
rect 324648 279460 324654 279472
rect 511258 279460 511264 279472
rect 324648 279432 511264 279460
rect 324648 279420 324654 279432
rect 511258 279420 511264 279432
rect 511316 279420 511322 279472
rect 317598 278128 317604 278180
rect 317656 278168 317662 278180
rect 477494 278168 477500 278180
rect 317656 278140 477500 278168
rect 317656 278128 317662 278140
rect 477494 278128 477500 278140
rect 477552 278128 477558 278180
rect 323210 278060 323216 278112
rect 323268 278100 323274 278112
rect 509234 278100 509240 278112
rect 323268 278072 509240 278100
rect 323268 278060 323274 278072
rect 509234 278060 509240 278072
rect 509292 278060 509298 278112
rect 35158 277992 35164 278044
rect 35216 278032 35222 278044
rect 236086 278032 236092 278044
rect 35216 278004 236092 278032
rect 35216 277992 35222 278004
rect 236086 277992 236092 278004
rect 236144 277992 236150 278044
rect 330386 277992 330392 278044
rect 330444 278032 330450 278044
rect 542354 278032 542360 278044
rect 330444 278004 542360 278032
rect 330444 277992 330450 278004
rect 542354 277992 542360 278004
rect 542412 277992 542418 278044
rect 310790 276700 310796 276752
rect 310848 276740 310854 276752
rect 440234 276740 440240 276752
rect 310848 276712 440240 276740
rect 310848 276700 310854 276712
rect 440234 276700 440240 276712
rect 440292 276700 440298 276752
rect 35894 276632 35900 276684
rect 35952 276672 35958 276684
rect 236362 276672 236368 276684
rect 35952 276644 236368 276672
rect 35952 276632 35958 276644
rect 236362 276632 236368 276644
rect 236420 276632 236426 276684
rect 320450 276632 320456 276684
rect 320508 276672 320514 276684
rect 496078 276672 496084 276684
rect 320508 276644 496084 276672
rect 320508 276632 320514 276644
rect 496078 276632 496084 276644
rect 496136 276632 496142 276684
rect 310698 275408 310704 275460
rect 310756 275448 310762 275460
rect 444374 275448 444380 275460
rect 310756 275420 444380 275448
rect 310756 275408 310762 275420
rect 444374 275408 444380 275420
rect 444432 275408 444438 275460
rect 44174 275340 44180 275392
rect 44232 275380 44238 275392
rect 236730 275380 236736 275392
rect 44232 275352 236736 275380
rect 44232 275340 44238 275352
rect 236730 275340 236736 275352
rect 236788 275340 236794 275392
rect 321738 275340 321744 275392
rect 321796 275380 321802 275392
rect 499574 275380 499580 275392
rect 321796 275352 499580 275380
rect 321796 275340 321802 275352
rect 499574 275340 499580 275352
rect 499632 275340 499638 275392
rect 22738 275272 22744 275324
rect 22796 275312 22802 275324
rect 233510 275312 233516 275324
rect 22796 275284 233516 275312
rect 22796 275272 22802 275284
rect 233510 275272 233516 275284
rect 233568 275272 233574 275324
rect 327350 275272 327356 275324
rect 327408 275312 327414 275324
rect 531314 275312 531320 275324
rect 327408 275284 531320 275312
rect 327408 275272 327414 275284
rect 531314 275272 531320 275284
rect 531372 275272 531378 275324
rect 312078 274116 312084 274168
rect 312136 274156 312142 274168
rect 448606 274156 448612 274168
rect 312136 274128 448612 274156
rect 312136 274116 312142 274128
rect 448606 274116 448612 274128
rect 448664 274116 448670 274168
rect 323118 274048 323124 274100
rect 323176 274088 323182 274100
rect 506474 274088 506480 274100
rect 323176 274060 506480 274088
rect 323176 274048 323182 274060
rect 506474 274048 506480 274060
rect 506532 274048 506538 274100
rect 14458 273980 14464 274032
rect 14516 274020 14522 274032
rect 230934 274020 230940 274032
rect 14516 273992 230940 274020
rect 14516 273980 14522 273992
rect 230934 273980 230940 273992
rect 230992 273980 230998 274032
rect 328638 273980 328644 274032
rect 328696 274020 328702 274032
rect 536098 274020 536104 274032
rect 328696 273992 536104 274020
rect 328696 273980 328702 273992
rect 536098 273980 536104 273992
rect 536156 273980 536162 274032
rect 99282 273912 99288 273964
rect 99340 273952 99346 273964
rect 336826 273952 336832 273964
rect 99340 273924 336832 273952
rect 99340 273912 99346 273924
rect 336826 273912 336832 273924
rect 336884 273912 336890 273964
rect 367738 273164 367744 273216
rect 367796 273204 367802 273216
rect 579890 273204 579896 273216
rect 367796 273176 579896 273204
rect 367796 273164 367802 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 326154 272552 326160 272604
rect 326212 272592 326218 272604
rect 521654 272592 521660 272604
rect 326212 272564 521660 272592
rect 326212 272552 326218 272564
rect 521654 272552 521660 272564
rect 521712 272552 521718 272604
rect 50338 272484 50344 272536
rect 50396 272524 50402 272536
rect 238938 272524 238944 272536
rect 50396 272496 238944 272524
rect 50396 272484 50402 272496
rect 238938 272484 238944 272496
rect 238996 272484 239002 272536
rect 332778 272484 332784 272536
rect 332836 272524 332842 272536
rect 560938 272524 560944 272536
rect 332836 272496 560944 272524
rect 332836 272484 332842 272496
rect 560938 272484 560944 272496
rect 560996 272484 561002 272536
rect 311986 271192 311992 271244
rect 312044 271232 312050 271244
rect 450538 271232 450544 271244
rect 312044 271204 450544 271232
rect 312044 271192 312050 271204
rect 450538 271192 450544 271204
rect 450596 271192 450602 271244
rect 52454 271124 52460 271176
rect 52512 271164 52518 271176
rect 239306 271164 239312 271176
rect 52512 271136 239312 271164
rect 52512 271124 52518 271136
rect 239306 271124 239312 271136
rect 239364 271124 239370 271176
rect 328546 271124 328552 271176
rect 328604 271164 328610 271176
rect 540238 271164 540244 271176
rect 328604 271136 540244 271164
rect 328604 271124 328610 271136
rect 540238 271124 540244 271136
rect 540296 271124 540302 271176
rect 313458 269900 313464 269952
rect 313516 269940 313522 269952
rect 458174 269940 458180 269952
rect 313516 269912 458180 269940
rect 313516 269900 313522 269912
rect 458174 269900 458180 269912
rect 458232 269900 458238 269952
rect 327258 269832 327264 269884
rect 327316 269872 327322 269884
rect 528554 269872 528560 269884
rect 327316 269844 528560 269872
rect 327316 269832 327322 269844
rect 528554 269832 528560 269844
rect 528612 269832 528618 269884
rect 57330 269764 57336 269816
rect 57388 269804 57394 269816
rect 240226 269804 240232 269816
rect 57388 269776 240232 269804
rect 57388 269764 57394 269776
rect 240226 269764 240232 269776
rect 240284 269764 240290 269816
rect 331490 269764 331496 269816
rect 331548 269804 331554 269816
rect 552014 269804 552020 269816
rect 331548 269776 552020 269804
rect 331548 269764 331554 269776
rect 552014 269764 552020 269776
rect 552072 269764 552078 269816
rect 314930 268472 314936 268524
rect 314988 268512 314994 268524
rect 464338 268512 464344 268524
rect 314988 268484 464344 268512
rect 314988 268472 314994 268484
rect 464338 268472 464344 268484
rect 464396 268472 464402 268524
rect 328454 268404 328460 268456
rect 328512 268444 328518 268456
rect 539686 268444 539692 268456
rect 328512 268416 539692 268444
rect 328512 268404 328518 268416
rect 539686 268404 539692 268416
rect 539744 268404 539750 268456
rect 59354 268336 59360 268388
rect 59412 268376 59418 268388
rect 240502 268376 240508 268388
rect 59412 268348 240508 268376
rect 59412 268336 59418 268348
rect 240502 268336 240508 268348
rect 240560 268336 240566 268388
rect 331398 268336 331404 268388
rect 331456 268376 331462 268388
rect 556246 268376 556252 268388
rect 331456 268348 556252 268376
rect 331456 268336 331462 268348
rect 556246 268336 556252 268348
rect 556304 268336 556310 268388
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 224218 267696 224224 267708
rect 3016 267668 224224 267696
rect 3016 267656 3022 267668
rect 224218 267656 224224 267668
rect 224276 267656 224282 267708
rect 238294 267112 238300 267164
rect 238352 267152 238358 267164
rect 350810 267152 350816 267164
rect 238352 267124 350816 267152
rect 238352 267112 238358 267124
rect 350810 267112 350816 267124
rect 350868 267112 350874 267164
rect 317506 267044 317512 267096
rect 317564 267084 317570 267096
rect 476114 267084 476120 267096
rect 317564 267056 476120 267084
rect 317564 267044 317570 267056
rect 476114 267044 476120 267056
rect 476172 267044 476178 267096
rect 332686 266976 332692 267028
rect 332744 267016 332750 267028
rect 558914 267016 558920 267028
rect 332744 266988 558920 267016
rect 332744 266976 332750 266988
rect 558914 266976 558920 266988
rect 558972 266976 558978 267028
rect 318886 265752 318892 265804
rect 318944 265792 318950 265804
rect 488534 265792 488540 265804
rect 318944 265764 488540 265792
rect 318944 265752 318950 265764
rect 488534 265752 488540 265764
rect 488592 265752 488598 265804
rect 331306 265684 331312 265736
rect 331364 265724 331370 265736
rect 554038 265724 554044 265736
rect 331364 265696 554044 265724
rect 331364 265684 331370 265696
rect 554038 265684 554044 265696
rect 554096 265684 554102 265736
rect 62114 265616 62120 265668
rect 62172 265656 62178 265668
rect 241606 265656 241612 265668
rect 62172 265628 241612 265656
rect 62172 265616 62178 265628
rect 241606 265616 241612 265628
rect 241664 265616 241670 265668
rect 335722 265616 335728 265668
rect 335780 265656 335786 265668
rect 574738 265656 574744 265668
rect 335780 265628 574744 265656
rect 335780 265616 335786 265628
rect 574738 265616 574744 265628
rect 574796 265616 574802 265668
rect 309594 264392 309600 264444
rect 309652 264432 309658 264444
rect 436738 264432 436744 264444
rect 309652 264404 436744 264432
rect 309652 264392 309658 264404
rect 436738 264392 436744 264404
rect 436796 264392 436802 264444
rect 310606 264324 310612 264376
rect 310664 264364 310670 264376
rect 440326 264364 440332 264376
rect 310664 264336 440332 264364
rect 310664 264324 310670 264336
rect 440326 264324 440332 264336
rect 440384 264324 440390 264376
rect 314838 264256 314844 264308
rect 314896 264296 314902 264308
rect 463694 264296 463700 264308
rect 314896 264268 463700 264296
rect 314896 264256 314902 264268
rect 463694 264256 463700 264268
rect 463752 264256 463758 264308
rect 66254 264188 66260 264240
rect 66312 264228 66318 264240
rect 241882 264228 241888 264240
rect 66312 264200 241888 264228
rect 66312 264188 66318 264200
rect 241882 264188 241888 264200
rect 241940 264188 241946 264240
rect 320358 264188 320364 264240
rect 320416 264228 320422 264240
rect 491294 264228 491300 264240
rect 320416 264200 491300 264228
rect 320416 264188 320422 264200
rect 491294 264188 491300 264200
rect 491352 264188 491358 264240
rect 238386 263032 238392 263084
rect 238444 263072 238450 263084
rect 360378 263072 360384 263084
rect 238444 263044 360384 263072
rect 238444 263032 238450 263044
rect 360378 263032 360384 263044
rect 360436 263032 360442 263084
rect 314746 262964 314752 263016
rect 314804 263004 314810 263016
rect 456058 263004 456064 263016
rect 314804 262976 456064 263004
rect 314804 262964 314810 262976
rect 456058 262964 456064 262976
rect 456116 262964 456122 263016
rect 75178 262896 75184 262948
rect 75236 262936 75242 262948
rect 243262 262936 243268 262948
rect 75236 262908 243268 262936
rect 75236 262896 75242 262908
rect 243262 262896 243268 262908
rect 243320 262896 243326 262948
rect 318794 262896 318800 262948
rect 318852 262936 318858 262948
rect 490006 262936 490012 262948
rect 318852 262908 490012 262936
rect 318852 262896 318858 262908
rect 490006 262896 490012 262908
rect 490064 262896 490070 262948
rect 4154 262828 4160 262880
rect 4212 262868 4218 262880
rect 229738 262868 229744 262880
rect 4212 262840 229744 262868
rect 4212 262828 4218 262840
rect 229738 262828 229744 262840
rect 229796 262828 229802 262880
rect 320266 262828 320272 262880
rect 320324 262868 320330 262880
rect 495434 262868 495440 262880
rect 320324 262840 495440 262868
rect 320324 262828 320330 262840
rect 495434 262828 495440 262840
rect 495492 262828 495498 262880
rect 320174 261604 320180 261656
rect 320232 261644 320238 261656
rect 492674 261644 492680 261656
rect 320232 261616 492680 261644
rect 320232 261604 320238 261616
rect 492674 261604 492680 261616
rect 492732 261604 492738 261656
rect 77294 261536 77300 261588
rect 77352 261576 77358 261588
rect 243170 261576 243176 261588
rect 77352 261548 243176 261576
rect 77352 261536 77358 261548
rect 243170 261536 243176 261548
rect 243228 261536 243234 261588
rect 321646 261536 321652 261588
rect 321704 261576 321710 261588
rect 494790 261576 494796 261588
rect 321704 261548 494796 261576
rect 321704 261536 321710 261548
rect 494790 261536 494796 261548
rect 494848 261536 494854 261588
rect 21358 261468 21364 261520
rect 21416 261508 21422 261520
rect 233418 261508 233424 261520
rect 21416 261480 233424 261508
rect 21416 261468 21422 261480
rect 233418 261468 233424 261480
rect 233476 261468 233482 261520
rect 330294 261468 330300 261520
rect 330352 261508 330358 261520
rect 546494 261508 546500 261520
rect 330352 261480 546500 261508
rect 330352 261468 330358 261480
rect 546494 261468 546500 261480
rect 546552 261468 546558 261520
rect 364978 260176 364984 260228
rect 365036 260216 365042 260228
rect 580442 260216 580448 260228
rect 365036 260188 580448 260216
rect 365036 260176 365042 260188
rect 580442 260176 580448 260188
rect 580500 260176 580506 260228
rect 42794 260108 42800 260160
rect 42852 260148 42858 260160
rect 237466 260148 237472 260160
rect 42852 260120 237472 260148
rect 42852 260108 42858 260120
rect 237466 260108 237472 260120
rect 237524 260108 237530 260160
rect 330202 260108 330208 260160
rect 330260 260148 330266 260160
rect 549254 260148 549260 260160
rect 330260 260120 549260 260148
rect 330260 260108 330266 260120
rect 549254 260108 549260 260120
rect 549312 260108 549318 260160
rect 91094 258748 91100 258800
rect 91152 258788 91158 258800
rect 246022 258788 246028 258800
rect 91152 258760 246028 258788
rect 91152 258748 91158 258760
rect 246022 258748 246028 258760
rect 246080 258748 246086 258800
rect 313366 258748 313372 258800
rect 313424 258788 313430 258800
rect 452654 258788 452660 258800
rect 313424 258760 452660 258788
rect 313424 258748 313430 258760
rect 452654 258748 452660 258760
rect 452712 258748 452718 258800
rect 13814 258680 13820 258732
rect 13872 258720 13878 258732
rect 231946 258720 231952 258732
rect 13872 258692 231952 258720
rect 13872 258680 13878 258692
rect 231946 258680 231952 258692
rect 232004 258680 232010 258732
rect 363598 258680 363604 258732
rect 363656 258720 363662 258732
rect 580350 258720 580356 258732
rect 363656 258692 580356 258720
rect 363656 258680 363662 258692
rect 580350 258680 580356 258692
rect 580408 258680 580414 258732
rect 326062 257388 326068 257440
rect 326120 257428 326126 257440
rect 527174 257428 527180 257440
rect 326120 257400 527180 257428
rect 326120 257388 326126 257400
rect 527174 257388 527180 257400
rect 527232 257388 527238 257440
rect 373258 257320 373264 257372
rect 373316 257360 373322 257372
rect 581086 257360 581092 257372
rect 373316 257332 581092 257360
rect 373316 257320 373322 257332
rect 581086 257320 581092 257332
rect 581144 257320 581150 257372
rect 325970 255960 325976 256012
rect 326028 256000 326034 256012
rect 523034 256000 523040 256012
rect 326028 255972 523040 256000
rect 326028 255960 326034 255972
rect 523034 255960 523040 255972
rect 523092 255960 523098 256012
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 220078 255252 220084 255264
rect 3200 255224 220084 255252
rect 3200 255212 3206 255224
rect 220078 255212 220084 255224
rect 220136 255212 220142 255264
rect 316034 254668 316040 254720
rect 316092 254708 316098 254720
rect 471974 254708 471980 254720
rect 316092 254680 471980 254708
rect 316092 254668 316098 254680
rect 471974 254668 471980 254680
rect 472032 254668 472038 254720
rect 317414 254600 317420 254652
rect 317472 254640 317478 254652
rect 478138 254640 478144 254652
rect 317472 254612 478144 254640
rect 317472 254600 317478 254612
rect 478138 254600 478144 254612
rect 478196 254600 478202 254652
rect 88334 254532 88340 254584
rect 88392 254572 88398 254584
rect 236638 254572 236644 254584
rect 88392 254544 236644 254572
rect 88392 254532 88398 254544
rect 236638 254532 236644 254544
rect 236696 254532 236702 254584
rect 330110 254532 330116 254584
rect 330168 254572 330174 254584
rect 547874 254572 547880 254584
rect 330168 254544 547880 254572
rect 330168 254532 330174 254544
rect 547874 254532 547880 254544
rect 547932 254532 547938 254584
rect 297726 253308 297732 253360
rect 297784 253348 297790 253360
rect 335630 253348 335636 253360
rect 297784 253320 335636 253348
rect 297784 253308 297790 253320
rect 335630 253308 335636 253320
rect 335688 253308 335694 253360
rect 97994 253240 98000 253292
rect 98052 253280 98058 253292
rect 247494 253280 247500 253292
rect 98052 253252 247500 253280
rect 98052 253240 98058 253252
rect 247494 253240 247500 253252
rect 247552 253240 247558 253292
rect 335446 253240 335452 253292
rect 335504 253280 335510 253292
rect 574094 253280 574100 253292
rect 335504 253252 574100 253280
rect 335504 253240 335510 253252
rect 574094 253240 574100 253252
rect 574152 253240 574158 253292
rect 30374 253172 30380 253224
rect 30432 253212 30438 253224
rect 234982 253212 234988 253224
rect 30432 253184 234988 253212
rect 30432 253172 30438 253184
rect 234982 253172 234988 253184
rect 235040 253172 235046 253224
rect 335538 253172 335544 253224
rect 335596 253212 335602 253224
rect 578234 253212 578240 253224
rect 335596 253184 578240 253212
rect 335596 253172 335602 253184
rect 578234 253172 578240 253184
rect 578292 253172 578298 253224
rect 297266 252016 297272 252068
rect 297324 252056 297330 252068
rect 344002 252056 344008 252068
rect 297324 252028 344008 252056
rect 297324 252016 297330 252028
rect 344002 252016 344008 252028
rect 344060 252016 344066 252068
rect 323026 251948 323032 252000
rect 323084 251988 323090 252000
rect 510614 251988 510620 252000
rect 323084 251960 510620 251988
rect 323084 251948 323090 251960
rect 510614 251948 510620 251960
rect 510672 251948 510678 252000
rect 324498 251880 324504 251932
rect 324556 251920 324562 251932
rect 514110 251920 514116 251932
rect 324556 251892 514116 251920
rect 324556 251880 324562 251892
rect 514110 251880 514116 251892
rect 514168 251880 514174 251932
rect 17954 251812 17960 251864
rect 18012 251852 18018 251864
rect 233326 251852 233332 251864
rect 18012 251824 233332 251852
rect 18012 251812 18018 251824
rect 233326 251812 233332 251824
rect 233384 251812 233390 251864
rect 332594 251812 332600 251864
rect 332652 251852 332658 251864
rect 564526 251852 564532 251864
rect 332652 251824 564532 251852
rect 332652 251812 332658 251824
rect 564526 251812 564532 251824
rect 564584 251812 564590 251864
rect 238478 250724 238484 250776
rect 238536 250764 238542 250776
rect 356330 250764 356336 250776
rect 238536 250736 356336 250764
rect 238536 250724 238542 250736
rect 356330 250724 356336 250736
rect 356388 250724 356394 250776
rect 359366 250724 359372 250776
rect 359424 250764 359430 250776
rect 441706 250764 441712 250776
rect 359424 250736 441712 250764
rect 359424 250724 359430 250736
rect 441706 250724 441712 250736
rect 441764 250724 441770 250776
rect 310514 250656 310520 250708
rect 310572 250696 310578 250708
rect 441614 250696 441620 250708
rect 310572 250668 441620 250696
rect 310572 250656 310578 250668
rect 441614 250656 441620 250668
rect 441672 250656 441678 250708
rect 311894 250588 311900 250640
rect 311952 250628 311958 250640
rect 445754 250628 445760 250640
rect 311952 250600 445760 250628
rect 311952 250588 311958 250600
rect 445754 250588 445760 250600
rect 445812 250588 445818 250640
rect 321554 250520 321560 250572
rect 321612 250560 321618 250572
rect 503714 250560 503720 250572
rect 321612 250532 503720 250560
rect 321612 250520 321618 250532
rect 503714 250520 503720 250532
rect 503772 250520 503778 250572
rect 22094 250452 22100 250504
rect 22152 250492 22158 250504
rect 233694 250492 233700 250504
rect 22152 250464 233700 250492
rect 22152 250452 22158 250464
rect 233694 250452 233700 250464
rect 233752 250452 233758 250504
rect 330018 250452 330024 250504
rect 330076 250492 330082 250504
rect 545114 250492 545120 250504
rect 330076 250464 545120 250492
rect 330076 250452 330082 250464
rect 545114 250452 545120 250464
rect 545172 250452 545178 250504
rect 313274 249160 313280 249212
rect 313332 249200 313338 249212
rect 456886 249200 456892 249212
rect 313332 249172 456892 249200
rect 313332 249160 313338 249172
rect 456886 249160 456892 249172
rect 456944 249160 456950 249212
rect 314654 249092 314660 249144
rect 314712 249132 314718 249144
rect 466454 249132 466460 249144
rect 314712 249104 466460 249132
rect 314712 249092 314718 249104
rect 466454 249092 466460 249104
rect 466512 249092 466518 249144
rect 12434 249024 12440 249076
rect 12492 249064 12498 249076
rect 232222 249064 232228 249076
rect 12492 249036 232228 249064
rect 12492 249024 12498 249036
rect 232222 249024 232228 249036
rect 232280 249024 232286 249076
rect 335354 249024 335360 249076
rect 335412 249064 335418 249076
rect 571978 249064 571984 249076
rect 335412 249036 571984 249064
rect 335412 249024 335418 249036
rect 571978 249024 571984 249036
rect 572036 249024 572042 249076
rect 298830 248344 298836 248396
rect 298888 248384 298894 248396
rect 347958 248384 347964 248396
rect 298888 248356 347964 248384
rect 298888 248344 298894 248356
rect 347958 248344 347964 248356
rect 348016 248344 348022 248396
rect 360286 248344 360292 248396
rect 360344 248384 360350 248396
rect 438210 248384 438216 248396
rect 360344 248356 438216 248384
rect 360344 248344 360350 248356
rect 438210 248344 438216 248356
rect 438268 248344 438274 248396
rect 292482 248276 292488 248328
rect 292540 248316 292546 248328
rect 345198 248316 345204 248328
rect 292540 248288 345204 248316
rect 292540 248276 292546 248288
rect 345198 248276 345204 248288
rect 345256 248276 345262 248328
rect 356238 248276 356244 248328
rect 356296 248316 356302 248328
rect 436922 248316 436928 248328
rect 356296 248288 436928 248316
rect 356296 248276 356302 248288
rect 436922 248276 436928 248288
rect 436980 248276 436986 248328
rect 297818 248208 297824 248260
rect 297876 248248 297882 248260
rect 350718 248248 350724 248260
rect 297876 248220 350724 248248
rect 297876 248208 297882 248220
rect 350718 248208 350724 248220
rect 350776 248208 350782 248260
rect 359274 248208 359280 248260
rect 359332 248248 359338 248260
rect 441798 248248 441804 248260
rect 359332 248220 441804 248248
rect 359332 248208 359338 248220
rect 441798 248208 441804 248220
rect 441856 248208 441862 248260
rect 286686 248140 286692 248192
rect 286744 248180 286750 248192
rect 346670 248180 346676 248192
rect 286744 248152 346676 248180
rect 286744 248140 286750 248152
rect 346670 248140 346676 248152
rect 346728 248140 346734 248192
rect 357802 248140 357808 248192
rect 357860 248180 357866 248192
rect 440602 248180 440608 248192
rect 357860 248152 440608 248180
rect 357860 248140 357866 248152
rect 440602 248140 440608 248152
rect 440660 248140 440666 248192
rect 288158 248072 288164 248124
rect 288216 248112 288222 248124
rect 348234 248112 348240 248124
rect 288216 248084 348240 248112
rect 288216 248072 288222 248084
rect 348234 248072 348240 248084
rect 348292 248072 348298 248124
rect 357710 248072 357716 248124
rect 357768 248112 357774 248124
rect 441890 248112 441896 248124
rect 357768 248084 441896 248112
rect 357768 248072 357774 248084
rect 441890 248072 441896 248084
rect 441948 248072 441954 248124
rect 288066 248004 288072 248056
rect 288124 248044 288130 248056
rect 305454 248044 305460 248056
rect 288124 248016 305460 248044
rect 288124 248004 288130 248016
rect 305454 248004 305460 248016
rect 305512 248004 305518 248056
rect 306926 248004 306932 248056
rect 306984 248044 306990 248056
rect 437474 248044 437480 248056
rect 306984 248016 437480 248044
rect 306984 248004 306990 248016
rect 437474 248004 437480 248016
rect 437532 248004 437538 248056
rect 289170 247936 289176 247988
rect 289228 247976 289234 247988
rect 303890 247976 303896 247988
rect 289228 247948 303896 247976
rect 289228 247936 289234 247948
rect 303890 247936 303896 247948
rect 303948 247936 303954 247988
rect 308214 247936 308220 247988
rect 308272 247976 308278 247988
rect 438854 247976 438860 247988
rect 308272 247948 438860 247976
rect 308272 247936 308278 247948
rect 438854 247936 438860 247948
rect 438912 247936 438918 247988
rect 290642 247868 290648 247920
rect 290700 247908 290706 247920
rect 305178 247908 305184 247920
rect 290700 247880 305184 247908
rect 290700 247868 290706 247880
rect 305178 247868 305184 247880
rect 305236 247868 305242 247920
rect 309502 247868 309508 247920
rect 309560 247908 309566 247920
rect 440418 247908 440424 247920
rect 309560 247880 440424 247908
rect 309560 247868 309566 247880
rect 440418 247868 440424 247880
rect 440476 247868 440482 247920
rect 292390 247800 292396 247852
rect 292448 247840 292454 247852
rect 305362 247840 305368 247852
rect 292448 247812 305368 247840
rect 292448 247800 292454 247812
rect 305362 247800 305368 247812
rect 305420 247800 305426 247852
rect 322934 247800 322940 247852
rect 322992 247840 322998 247852
rect 506566 247840 506572 247852
rect 322992 247812 506572 247840
rect 322992 247800 322998 247812
rect 506566 247800 506572 247812
rect 506624 247800 506630 247852
rect 324406 247732 324412 247784
rect 324464 247772 324470 247784
rect 517514 247772 517520 247784
rect 324464 247744 517520 247772
rect 324464 247732 324470 247744
rect 517514 247732 517520 247744
rect 517572 247732 517578 247784
rect 4798 247664 4804 247716
rect 4856 247704 4862 247716
rect 229186 247704 229192 247716
rect 4856 247676 229192 247704
rect 4856 247664 4862 247676
rect 229186 247664 229192 247676
rect 229244 247664 229250 247716
rect 287882 247664 287888 247716
rect 287940 247704 287946 247716
rect 300670 247704 300676 247716
rect 287940 247676 300676 247704
rect 287940 247664 287946 247676
rect 300670 247664 300676 247676
rect 300728 247664 300734 247716
rect 329926 247664 329932 247716
rect 329984 247704 329990 247716
rect 547966 247704 547972 247716
rect 329984 247676 547972 247704
rect 329984 247664 329990 247676
rect 547966 247664 547972 247676
rect 548024 247664 548030 247716
rect 300762 247596 300768 247648
rect 300820 247636 300826 247648
rect 346762 247636 346768 247648
rect 300820 247608 346768 247636
rect 300820 247596 300826 247608
rect 346762 247596 346768 247608
rect 346820 247596 346826 247648
rect 297082 247528 297088 247580
rect 297140 247568 297146 247580
rect 339586 247568 339592 247580
rect 297140 247540 339592 247568
rect 297140 247528 297146 247540
rect 339586 247528 339592 247540
rect 339644 247528 339650 247580
rect 288986 247460 288992 247512
rect 289044 247500 289050 247512
rect 303798 247500 303804 247512
rect 289044 247472 303804 247500
rect 289044 247460 289050 247472
rect 303798 247460 303804 247472
rect 303856 247460 303862 247512
rect 286778 247392 286784 247444
rect 286836 247432 286842 247444
rect 303982 247432 303988 247444
rect 286836 247404 303988 247432
rect 286836 247392 286842 247404
rect 303982 247392 303988 247404
rect 304040 247392 304046 247444
rect 298738 247052 298744 247104
rect 298796 247092 298802 247104
rect 304074 247092 304080 247104
rect 298796 247064 304080 247092
rect 298796 247052 298802 247064
rect 304074 247052 304080 247064
rect 304132 247052 304138 247104
rect 297358 246984 297364 247036
rect 297416 247024 297422 247036
rect 342714 247024 342720 247036
rect 297416 246996 342720 247024
rect 297416 246984 297422 246996
rect 342714 246984 342720 246996
rect 342772 246984 342778 247036
rect 298922 246916 298928 246968
rect 298980 246956 298986 246968
rect 345474 246956 345480 246968
rect 298980 246928 345480 246956
rect 298980 246916 298986 246928
rect 345474 246916 345480 246928
rect 345532 246916 345538 246968
rect 299382 246848 299388 246900
rect 299440 246888 299446 246900
rect 350994 246888 351000 246900
rect 299440 246860 351000 246888
rect 299440 246848 299446 246860
rect 350994 246848 351000 246860
rect 351052 246848 351058 246900
rect 297174 246780 297180 246832
rect 297232 246820 297238 246832
rect 349430 246820 349436 246832
rect 297232 246792 349436 246820
rect 297232 246780 297238 246792
rect 349430 246780 349436 246792
rect 349488 246780 349494 246832
rect 296530 246712 296536 246764
rect 296588 246752 296594 246764
rect 350902 246752 350908 246764
rect 296588 246724 350908 246752
rect 296588 246712 296594 246724
rect 350902 246712 350908 246724
rect 350960 246712 350966 246764
rect 289630 246644 289636 246696
rect 289688 246684 289694 246696
rect 349246 246684 349252 246696
rect 289688 246656 349252 246684
rect 289688 246644 289694 246656
rect 349246 246644 349252 246656
rect 349304 246644 349310 246696
rect 325878 246576 325884 246628
rect 325936 246616 325942 246628
rect 524414 246616 524420 246628
rect 325936 246588 524420 246616
rect 325936 246576 325942 246588
rect 524414 246576 524420 246588
rect 524472 246576 524478 246628
rect 325786 246508 325792 246560
rect 325844 246548 325850 246560
rect 525794 246548 525800 246560
rect 325844 246520 525800 246548
rect 325844 246508 325850 246520
rect 525794 246508 525800 246520
rect 525852 246508 525858 246560
rect 327166 246440 327172 246492
rect 327224 246480 327230 246492
rect 534074 246480 534080 246492
rect 327224 246452 534080 246480
rect 327224 246440 327230 246452
rect 534074 246440 534080 246452
rect 534132 246440 534138 246492
rect 329834 246372 329840 246424
rect 329892 246412 329898 246424
rect 543734 246412 543740 246424
rect 329892 246384 543740 246412
rect 329892 246372 329898 246384
rect 543734 246372 543740 246384
rect 543792 246372 543798 246424
rect 3602 246304 3608 246356
rect 3660 246344 3666 246356
rect 228358 246344 228364 246356
rect 3660 246316 228364 246344
rect 3660 246304 3666 246316
rect 228358 246304 228364 246316
rect 228416 246304 228422 246356
rect 331214 246304 331220 246356
rect 331272 246344 331278 246356
rect 553394 246344 553400 246356
rect 331272 246316 553400 246344
rect 331272 246304 331278 246316
rect 553394 246304 553400 246316
rect 553452 246304 553458 246356
rect 297450 246236 297456 246288
rect 297508 246276 297514 246288
rect 341150 246276 341156 246288
rect 297508 246248 341156 246276
rect 297508 246236 297514 246248
rect 341150 246236 341156 246248
rect 341208 246236 341214 246288
rect 291010 245556 291016 245608
rect 291068 245596 291074 245608
rect 306650 245596 306656 245608
rect 291068 245568 306656 245596
rect 291068 245556 291074 245568
rect 306650 245556 306656 245568
rect 306708 245556 306714 245608
rect 309410 245556 309416 245608
rect 309468 245596 309474 245608
rect 437934 245596 437940 245608
rect 309468 245568 437940 245596
rect 309468 245556 309474 245568
rect 437934 245556 437940 245568
rect 437992 245556 437998 245608
rect 292206 245488 292212 245540
rect 292264 245528 292270 245540
rect 305086 245528 305092 245540
rect 292264 245500 305092 245528
rect 292264 245488 292270 245500
rect 305086 245488 305092 245500
rect 305144 245488 305150 245540
rect 307938 245488 307944 245540
rect 307996 245528 308002 245540
rect 437658 245528 437664 245540
rect 307996 245500 437664 245528
rect 307996 245488 308002 245500
rect 437658 245488 437664 245500
rect 437716 245488 437722 245540
rect 293678 245420 293684 245472
rect 293736 245460 293742 245472
rect 303706 245460 303712 245472
rect 293736 245432 303712 245460
rect 293736 245420 293742 245432
rect 303706 245420 303712 245432
rect 303764 245420 303770 245472
rect 309318 245420 309324 245472
rect 309376 245460 309382 245472
rect 439130 245460 439136 245472
rect 309376 245432 439136 245460
rect 309376 245420 309382 245432
rect 439130 245420 439136 245432
rect 439188 245420 439194 245472
rect 293402 245352 293408 245404
rect 293460 245392 293466 245404
rect 303614 245392 303620 245404
rect 293460 245364 303620 245392
rect 293460 245352 293466 245364
rect 303614 245352 303620 245364
rect 303672 245352 303678 245404
rect 307846 245352 307852 245404
rect 307904 245392 307910 245404
rect 437842 245392 437848 245404
rect 307904 245364 437848 245392
rect 307904 245352 307910 245364
rect 437842 245352 437848 245364
rect 437900 245352 437906 245404
rect 295242 245284 295248 245336
rect 295300 245324 295306 245336
rect 304994 245324 305000 245336
rect 295300 245296 305000 245324
rect 295300 245284 295306 245296
rect 304994 245284 305000 245296
rect 305052 245284 305058 245336
rect 309134 245284 309140 245336
rect 309192 245324 309198 245336
rect 439314 245324 439320 245336
rect 309192 245296 439320 245324
rect 309192 245284 309198 245296
rect 439314 245284 439320 245296
rect 439372 245284 439378 245336
rect 306834 245216 306840 245268
rect 306892 245256 306898 245268
rect 437566 245256 437572 245268
rect 306892 245228 437572 245256
rect 306892 245216 306898 245228
rect 437566 245216 437572 245228
rect 437624 245216 437630 245268
rect 295150 245148 295156 245200
rect 295208 245188 295214 245200
rect 300854 245188 300860 245200
rect 295208 245160 300860 245188
rect 295208 245148 295214 245160
rect 300854 245148 300860 245160
rect 300912 245148 300918 245200
rect 306466 245148 306472 245200
rect 306524 245188 306530 245200
rect 437750 245188 437756 245200
rect 306524 245160 437756 245188
rect 306524 245148 306530 245160
rect 437750 245148 437756 245160
rect 437808 245148 437814 245200
rect 292482 245080 292488 245132
rect 292540 245120 292546 245132
rect 299566 245120 299572 245132
rect 292540 245092 299572 245120
rect 292540 245080 292546 245092
rect 299566 245080 299572 245092
rect 299624 245080 299630 245132
rect 308030 245080 308036 245132
rect 308088 245120 308094 245132
rect 439406 245120 439412 245132
rect 308088 245092 439412 245120
rect 308088 245080 308094 245092
rect 439406 245080 439412 245092
rect 439464 245080 439470 245132
rect 291102 245012 291108 245064
rect 291160 245052 291166 245064
rect 299658 245052 299664 245064
rect 291160 245024 299664 245052
rect 291160 245012 291166 245024
rect 299658 245012 299664 245024
rect 299716 245012 299722 245064
rect 307754 245012 307760 245064
rect 307812 245052 307818 245064
rect 439222 245052 439228 245064
rect 307812 245024 439228 245052
rect 307812 245012 307818 245024
rect 439222 245012 439228 245024
rect 439280 245012 439286 245064
rect 291010 244944 291016 244996
rect 291068 244984 291074 244996
rect 301130 244984 301136 244996
rect 291068 244956 301136 244984
rect 291068 244944 291074 244956
rect 301130 244944 301136 244956
rect 301188 244944 301194 244996
rect 306742 244944 306748 244996
rect 306800 244984 306806 244996
rect 438946 244984 438952 244996
rect 306800 244956 438952 244984
rect 306800 244944 306806 244956
rect 438946 244944 438952 244956
rect 439004 244944 439010 244996
rect 7650 244876 7656 244928
rect 7708 244916 7714 244928
rect 230842 244916 230848 244928
rect 7708 244888 230848 244916
rect 7708 244876 7714 244888
rect 230842 244876 230848 244888
rect 230900 244876 230906 244928
rect 289722 244876 289728 244928
rect 289780 244916 289786 244928
rect 302234 244916 302240 244928
rect 289780 244888 302240 244916
rect 289780 244876 289786 244888
rect 302234 244876 302240 244888
rect 302292 244876 302298 244928
rect 306374 244876 306380 244928
rect 306432 244916 306438 244928
rect 439038 244916 439044 244928
rect 306432 244888 439044 244916
rect 306432 244876 306438 244888
rect 439038 244876 439044 244888
rect 439096 244876 439102 244928
rect 299106 244808 299112 244860
rect 299164 244848 299170 244860
rect 342622 244848 342628 244860
rect 299164 244820 342628 244848
rect 299164 244808 299170 244820
rect 342622 244808 342628 244820
rect 342680 244808 342686 244860
rect 356514 244808 356520 244860
rect 356572 244848 356578 244860
rect 438302 244848 438308 244860
rect 356572 244820 438308 244848
rect 356572 244808 356578 244820
rect 438302 244808 438308 244820
rect 438360 244808 438366 244860
rect 299014 244740 299020 244792
rect 299072 244780 299078 244792
rect 339770 244780 339776 244792
rect 299072 244752 339776 244780
rect 299072 244740 299078 244752
rect 339770 244740 339776 244752
rect 339828 244740 339834 244792
rect 360470 244740 360476 244792
rect 360528 244780 360534 244792
rect 439682 244780 439688 244792
rect 360528 244752 439688 244780
rect 360528 244740 360534 244752
rect 439682 244740 439688 244752
rect 439740 244740 439746 244792
rect 297634 244672 297640 244724
rect 297692 244712 297698 244724
rect 337010 244712 337016 244724
rect 297692 244684 337016 244712
rect 297692 244672 297698 244684
rect 337010 244672 337016 244684
rect 337068 244672 337074 244724
rect 295242 244604 295248 244656
rect 295300 244644 295306 244656
rect 299474 244644 299480 244656
rect 295300 244616 299480 244644
rect 295300 244604 295306 244616
rect 299474 244604 299480 244616
rect 299532 244604 299538 244656
rect 288342 244468 288348 244520
rect 288400 244508 288406 244520
rect 291746 244508 291752 244520
rect 288400 244480 291752 244508
rect 288400 244468 288406 244480
rect 291746 244468 291752 244480
rect 291804 244468 291810 244520
rect 291746 244332 291752 244384
rect 291804 244372 291810 244384
rect 299290 244372 299296 244384
rect 291804 244344 299296 244372
rect 291804 244332 291810 244344
rect 299290 244332 299296 244344
rect 299348 244332 299354 244384
rect 293678 243720 293684 243772
rect 293736 243760 293742 243772
rect 300762 243760 300768 243772
rect 293736 243732 300768 243760
rect 293736 243720 293742 243732
rect 300762 243720 300768 243732
rect 300820 243720 300826 243772
rect 299290 243652 299296 243704
rect 299348 243692 299354 243704
rect 343910 243692 343916 243704
rect 299348 243664 343916 243692
rect 299348 243652 299354 243664
rect 343910 243652 343916 243664
rect 343968 243652 343974 243704
rect 299198 243584 299204 243636
rect 299256 243624 299262 243636
rect 345382 243624 345388 243636
rect 299256 243596 345388 243624
rect 299256 243584 299262 243596
rect 345382 243584 345388 243596
rect 345440 243584 345446 243636
rect 97810 243516 97816 243568
rect 97868 243556 97874 243568
rect 297266 243556 297272 243568
rect 97868 243528 297272 243556
rect 97868 243516 97874 243528
rect 297266 243516 297272 243528
rect 297324 243516 297330 243568
rect 297910 243516 297916 243568
rect 297968 243556 297974 243568
rect 356054 243556 356060 243568
rect 297968 243528 356060 243556
rect 297968 243516 297974 243528
rect 356054 243516 356060 243528
rect 356112 243516 356118 243568
rect 97902 243448 97908 243500
rect 97960 243488 97966 243500
rect 298738 243488 298744 243500
rect 97960 243460 298744 243488
rect 97960 243448 97966 243460
rect 298738 243448 298744 243460
rect 298796 243488 298802 243500
rect 299014 243488 299020 243500
rect 298796 243460 299020 243488
rect 298796 243448 298802 243460
rect 299014 243448 299020 243460
rect 299072 243448 299078 243500
rect 97718 243380 97724 243432
rect 97776 243420 97782 243432
rect 298922 243420 298928 243432
rect 97776 243392 298928 243420
rect 97776 243380 97782 243392
rect 298922 243380 298928 243392
rect 298980 243380 298986 243432
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 98638 241448 98644 241460
rect 3292 241420 98644 241448
rect 3292 241408 3298 241420
rect 98638 241408 98644 241420
rect 98696 241408 98702 241460
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 86218 215268 86224 215280
rect 3384 215240 86224 215268
rect 3384 215228 3390 215240
rect 86218 215228 86224 215240
rect 86276 215228 86282 215280
rect 292206 198024 292212 198076
rect 292264 198064 292270 198076
rect 297174 198064 297180 198076
rect 292264 198036 297180 198064
rect 292264 198024 292270 198036
rect 297174 198024 297180 198036
rect 297232 198024 297238 198076
rect 297542 197412 297548 197464
rect 297600 197452 297606 197464
rect 298830 197452 298836 197464
rect 297600 197424 298836 197452
rect 297600 197412 297606 197424
rect 298830 197412 298836 197424
rect 298888 197412 298894 197464
rect 292390 197276 292396 197328
rect 292448 197316 292454 197328
rect 298830 197316 298836 197328
rect 292448 197288 298836 197316
rect 292448 197276 292454 197288
rect 298830 197276 298836 197288
rect 298888 197276 298894 197328
rect 296622 195916 296628 195968
rect 296680 195956 296686 195968
rect 298370 195956 298376 195968
rect 296680 195928 298376 195956
rect 296680 195916 296686 195928
rect 298370 195916 298376 195928
rect 298428 195916 298434 195968
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 95970 189020 95976 189032
rect 3200 188992 95976 189020
rect 3200 188980 3206 188992
rect 95970 188980 95976 188992
rect 96028 188980 96034 189032
rect 261110 177284 261116 177336
rect 261168 177324 261174 177336
rect 277670 177324 277676 177336
rect 261168 177296 277676 177324
rect 261168 177284 261174 177296
rect 277670 177284 277676 177296
rect 277728 177284 277734 177336
rect 285214 171028 285220 171080
rect 285272 171068 285278 171080
rect 297174 171068 297180 171080
rect 285272 171040 297180 171068
rect 285272 171028 285278 171040
rect 297174 171028 297180 171040
rect 297232 171028 297238 171080
rect 236730 170348 236736 170400
rect 236788 170388 236794 170400
rect 285214 170388 285220 170400
rect 236788 170360 285220 170388
rect 236788 170348 236794 170360
rect 285214 170348 285220 170360
rect 285272 170348 285278 170400
rect 238570 167628 238576 167680
rect 238628 167668 238634 167680
rect 297726 167668 297732 167680
rect 238628 167640 297732 167668
rect 238628 167628 238634 167640
rect 297726 167628 297732 167640
rect 297784 167628 297790 167680
rect 292298 166948 292304 167000
rect 292356 166988 292362 167000
rect 296714 166988 296720 167000
rect 292356 166960 296720 166988
rect 292356 166948 292362 166960
rect 296714 166948 296720 166960
rect 296772 166948 296778 167000
rect 3510 164160 3516 164212
rect 3568 164200 3574 164212
rect 84838 164200 84844 164212
rect 3568 164172 84844 164200
rect 3568 164160 3574 164172
rect 84838 164160 84844 164172
rect 84896 164160 84902 164212
rect 97810 159876 97816 159928
rect 97868 159916 97874 159928
rect 298922 159916 298928 159928
rect 97868 159888 298928 159916
rect 97868 159876 97874 159888
rect 298922 159876 298928 159888
rect 298980 159876 298986 159928
rect 97626 159808 97632 159860
rect 97684 159848 97690 159860
rect 297266 159848 297272 159860
rect 97684 159820 297272 159848
rect 97684 159808 97690 159820
rect 297266 159808 297272 159820
rect 297324 159808 297330 159860
rect 97534 159740 97540 159792
rect 97592 159780 97598 159792
rect 297358 159780 297364 159792
rect 97592 159752 297364 159780
rect 97592 159740 97598 159752
rect 297358 159740 297364 159752
rect 297416 159740 297422 159792
rect 97442 159672 97448 159724
rect 97500 159712 97506 159724
rect 238570 159712 238576 159724
rect 97500 159684 238576 159712
rect 97500 159672 97506 159684
rect 238570 159672 238576 159684
rect 238628 159672 238634 159724
rect 97902 159604 97908 159656
rect 97960 159644 97966 159656
rect 236730 159644 236736 159656
rect 97960 159616 236736 159644
rect 97960 159604 97966 159616
rect 236730 159604 236736 159616
rect 236788 159604 236794 159656
rect 284478 159604 284484 159656
rect 284536 159644 284542 159656
rect 299474 159644 299480 159656
rect 284536 159616 299480 159644
rect 284536 159604 284542 159616
rect 299474 159604 299480 159616
rect 299532 159604 299538 159656
rect 287606 159536 287612 159588
rect 287664 159576 287670 159588
rect 309134 159576 309140 159588
rect 287664 159548 309140 159576
rect 287664 159536 287670 159548
rect 309134 159536 309140 159548
rect 309192 159536 309198 159588
rect 293310 159468 293316 159520
rect 293368 159508 293374 159520
rect 327166 159508 327172 159520
rect 293368 159480 327172 159508
rect 293368 159468 293374 159480
rect 327166 159468 327172 159480
rect 327224 159468 327230 159520
rect 234614 159400 234620 159452
rect 234672 159440 234678 159452
rect 273714 159440 273720 159452
rect 234672 159412 273720 159440
rect 234672 159400 234678 159412
rect 273714 159400 273720 159412
rect 273772 159400 273778 159452
rect 298186 159400 298192 159452
rect 298244 159440 298250 159452
rect 338758 159440 338764 159452
rect 298244 159412 338764 159440
rect 298244 159400 298250 159412
rect 338758 159400 338764 159412
rect 338816 159400 338822 159452
rect 220814 159332 220820 159384
rect 220872 159372 220878 159384
rect 271046 159372 271052 159384
rect 220872 159344 271052 159372
rect 220872 159332 220878 159344
rect 271046 159332 271052 159344
rect 271104 159332 271110 159384
rect 298830 159332 298836 159384
rect 298888 159372 298894 159384
rect 348234 159372 348240 159384
rect 298888 159344 348240 159372
rect 298888 159332 298894 159344
rect 348234 159332 348240 159344
rect 348292 159332 348298 159384
rect 293678 159264 293684 159316
rect 293736 159304 293742 159316
rect 350994 159304 351000 159316
rect 293736 159276 351000 159304
rect 293736 159264 293742 159276
rect 350994 159264 351000 159276
rect 351052 159264 351058 159316
rect 297542 159196 297548 159248
rect 297600 159236 297606 159248
rect 356054 159236 356060 159248
rect 297600 159208 356060 159236
rect 297600 159196 297606 159208
rect 356054 159196 356060 159208
rect 356112 159196 356118 159248
rect 286778 159128 286784 159180
rect 286836 159168 286842 159180
rect 353570 159168 353576 159180
rect 286836 159140 353576 159168
rect 286836 159128 286842 159140
rect 353570 159128 353576 159140
rect 353628 159128 353634 159180
rect 165982 159060 165988 159112
rect 166040 159100 166046 159112
rect 238110 159100 238116 159112
rect 166040 159072 238116 159100
rect 166040 159060 166046 159072
rect 238110 159060 238116 159072
rect 238168 159060 238174 159112
rect 299382 159060 299388 159112
rect 299440 159100 299446 159112
rect 368290 159100 368296 159112
rect 299440 159072 368296 159100
rect 299440 159060 299446 159072
rect 368290 159060 368296 159072
rect 368348 159060 368354 159112
rect 160922 158992 160928 159044
rect 160980 159032 160986 159044
rect 240778 159032 240784 159044
rect 160980 159004 240784 159032
rect 160980 158992 160986 159004
rect 240778 158992 240784 159004
rect 240836 158992 240842 159044
rect 296530 158992 296536 159044
rect 296588 159032 296594 159044
rect 365898 159032 365904 159044
rect 296588 159004 365904 159032
rect 296588 158992 296594 159004
rect 365898 158992 365904 159004
rect 365956 158992 365962 159044
rect 156046 158924 156052 158976
rect 156104 158964 156110 158976
rect 249058 158964 249064 158976
rect 156104 158936 249064 158964
rect 156104 158924 156110 158936
rect 249058 158924 249064 158936
rect 249116 158924 249122 158976
rect 288158 158924 288164 158976
rect 288216 158964 288222 158976
rect 358446 158964 358452 158976
rect 288216 158936 358452 158964
rect 288216 158924 288222 158936
rect 358446 158924 358452 158936
rect 358504 158924 358510 158976
rect 153654 158856 153660 158908
rect 153712 158896 153718 158908
rect 250530 158896 250536 158908
rect 153712 158868 250536 158896
rect 153712 158856 153718 158868
rect 250530 158856 250536 158868
rect 250588 158856 250594 158908
rect 289630 158856 289636 158908
rect 289688 158896 289694 158908
rect 360930 158896 360936 158908
rect 289688 158868 360936 158896
rect 289688 158856 289694 158868
rect 360930 158856 360936 158868
rect 360988 158856 360994 158908
rect 168282 158788 168288 158840
rect 168340 158828 168346 158840
rect 286410 158828 286416 158840
rect 168340 158800 286416 158828
rect 168340 158788 168346 158800
rect 286410 158788 286416 158800
rect 286468 158788 286474 158840
rect 292206 158788 292212 158840
rect 292264 158828 292270 158840
rect 363414 158828 363420 158840
rect 292264 158800 363420 158828
rect 292264 158788 292270 158800
rect 363414 158788 363420 158800
rect 363472 158788 363478 158840
rect 175918 158720 175924 158772
rect 175976 158760 175982 158772
rect 296162 158760 296168 158772
rect 175976 158732 296168 158760
rect 175976 158720 175982 158732
rect 296162 158720 296168 158732
rect 296220 158720 296226 158772
rect 297818 158720 297824 158772
rect 297876 158760 297882 158772
rect 370958 158760 370964 158772
rect 297876 158732 370964 158760
rect 297876 158720 297882 158732
rect 370958 158720 370964 158732
rect 371016 158720 371022 158772
rect 388530 158720 388536 158772
rect 388588 158760 388594 158772
rect 436922 158760 436928 158772
rect 388588 158732 436928 158760
rect 388588 158720 388594 158732
rect 436922 158720 436928 158732
rect 436980 158720 436986 158772
rect 128722 158652 128728 158704
rect 128780 158692 128786 158704
rect 276014 158692 276020 158704
rect 128780 158664 276020 158692
rect 128780 158652 128786 158664
rect 276014 158652 276020 158664
rect 276072 158652 276078 158704
rect 293770 158652 293776 158704
rect 293828 158692 293834 158704
rect 338390 158692 338396 158704
rect 293828 158664 338396 158692
rect 293828 158652 293834 158664
rect 338390 158652 338396 158664
rect 338448 158652 338454 158704
rect 373442 158652 373448 158704
rect 373500 158692 373506 158704
rect 440510 158692 440516 158704
rect 373500 158664 440516 158692
rect 373500 158652 373506 158664
rect 440510 158652 440516 158664
rect 440568 158652 440574 158704
rect 126514 158584 126520 158636
rect 126572 158624 126578 158636
rect 276566 158624 276572 158636
rect 126572 158596 276572 158624
rect 126572 158584 126578 158596
rect 276566 158584 276572 158596
rect 276624 158624 276630 158636
rect 276842 158624 276848 158636
rect 276624 158596 276848 158624
rect 276624 158584 276630 158596
rect 276842 158584 276848 158596
rect 276900 158584 276906 158636
rect 298002 158584 298008 158636
rect 298060 158624 298066 158636
rect 331214 158624 331220 158636
rect 298060 158596 331220 158624
rect 298060 158584 298066 158596
rect 331214 158584 331220 158596
rect 331272 158584 331278 158636
rect 376018 158584 376024 158636
rect 376076 158624 376082 158636
rect 438118 158624 438124 158636
rect 376076 158596 438124 158624
rect 376076 158584 376082 158596
rect 438118 158584 438124 158596
rect 438176 158584 438182 158636
rect 121914 158516 121920 158568
rect 121972 158556 121978 158568
rect 290734 158556 290740 158568
rect 121972 158528 290740 158556
rect 121972 158516 121978 158528
rect 290734 158516 290740 158528
rect 290792 158516 290798 158568
rect 294966 158516 294972 158568
rect 295024 158556 295030 158568
rect 340966 158556 340972 158568
rect 295024 158528 340972 158556
rect 295024 158516 295030 158528
rect 340966 158516 340972 158528
rect 341024 158516 341030 158568
rect 378594 158516 378600 158568
rect 378652 158556 378658 158568
rect 439590 158556 439596 158568
rect 378652 158528 439596 158556
rect 378652 158516 378658 158528
rect 439590 158516 439596 158528
rect 439648 158516 439654 158568
rect 120626 158448 120632 158500
rect 120684 158488 120690 158500
rect 288250 158488 288256 158500
rect 120684 158460 288256 158488
rect 120684 158448 120690 158460
rect 288250 158448 288256 158460
rect 288308 158448 288314 158500
rect 290642 158448 290648 158500
rect 290700 158488 290706 158500
rect 290918 158488 290924 158500
rect 290700 158460 290924 158488
rect 290700 158448 290706 158460
rect 290918 158448 290924 158460
rect 290976 158448 290982 158500
rect 293586 158448 293592 158500
rect 293644 158488 293650 158500
rect 328270 158488 328276 158500
rect 293644 158460 328276 158488
rect 293644 158448 293650 158460
rect 328270 158448 328276 158460
rect 328328 158448 328334 158500
rect 380986 158448 380992 158500
rect 381044 158488 381050 158500
rect 436830 158488 436836 158500
rect 381044 158460 436836 158488
rect 381044 158448 381050 158460
rect 436830 158448 436836 158460
rect 436888 158448 436894 158500
rect 282454 158380 282460 158432
rect 282512 158420 282518 158432
rect 343542 158420 343548 158432
rect 282512 158392 343548 158420
rect 282512 158380 282518 158392
rect 343542 158380 343548 158392
rect 343600 158380 343606 158432
rect 383562 158380 383568 158432
rect 383620 158420 383626 158432
rect 438026 158420 438032 158432
rect 383620 158392 438032 158420
rect 383620 158380 383626 158392
rect 438026 158380 438032 158392
rect 438084 158380 438090 158432
rect 127618 158312 127624 158364
rect 127676 158352 127682 158364
rect 295058 158352 295064 158364
rect 127676 158324 295064 158352
rect 127676 158312 127682 158324
rect 295058 158312 295064 158324
rect 295116 158352 295122 158364
rect 327534 158352 327540 158364
rect 295116 158324 327540 158352
rect 295116 158312 295122 158324
rect 327534 158312 327540 158324
rect 327592 158312 327598 158364
rect 385954 158312 385960 158364
rect 386012 158352 386018 158364
rect 439498 158352 439504 158364
rect 386012 158324 439504 158352
rect 386012 158312 386018 158324
rect 439498 158312 439504 158324
rect 439556 158312 439562 158364
rect 132402 158244 132408 158296
rect 132460 158284 132466 158296
rect 299198 158284 299204 158296
rect 132460 158256 299204 158284
rect 132460 158244 132466 158256
rect 299198 158244 299204 158256
rect 299256 158284 299262 158296
rect 332318 158284 332324 158296
rect 299256 158256 332324 158284
rect 299256 158244 299262 158256
rect 332318 158244 332324 158256
rect 332376 158244 332382 158296
rect 391474 158244 391480 158296
rect 391532 158284 391538 158296
rect 438302 158284 438308 158296
rect 391532 158256 438308 158284
rect 391532 158244 391538 158256
rect 438302 158244 438308 158256
rect 438360 158244 438366 158296
rect 131298 158176 131304 158228
rect 131356 158216 131362 158228
rect 298002 158216 298008 158228
rect 131356 158188 298008 158216
rect 131356 158176 131362 158188
rect 298002 158176 298008 158188
rect 298060 158176 298066 158228
rect 299382 158176 299388 158228
rect 299440 158216 299446 158228
rect 329926 158216 329932 158228
rect 299440 158188 329932 158216
rect 299440 158176 299446 158188
rect 329926 158176 329932 158188
rect 329984 158176 329990 158228
rect 394234 158176 394240 158228
rect 394292 158216 394298 158228
rect 440602 158216 440608 158228
rect 394292 158188 440608 158216
rect 394292 158176 394298 158188
rect 440602 158176 440608 158188
rect 440660 158176 440666 158228
rect 275922 158108 275928 158160
rect 275980 158148 275986 158160
rect 335998 158148 336004 158160
rect 275980 158120 336004 158148
rect 275980 158108 275986 158120
rect 335998 158108 336004 158120
rect 336056 158108 336062 158160
rect 395890 158108 395896 158160
rect 395948 158148 395954 158160
rect 441890 158148 441896 158160
rect 395948 158120 441896 158148
rect 395948 158108 395954 158120
rect 441890 158108 441896 158120
rect 441948 158108 441954 158160
rect 133506 158040 133512 158092
rect 133564 158080 133570 158092
rect 283834 158080 283840 158092
rect 133564 158052 283840 158080
rect 133564 158040 133570 158052
rect 283834 158040 283840 158052
rect 283892 158040 283898 158092
rect 286134 158040 286140 158092
rect 286192 158080 286198 158092
rect 286870 158080 286876 158092
rect 286192 158052 286876 158080
rect 286192 158040 286198 158052
rect 286870 158040 286876 158052
rect 286928 158080 286934 158092
rect 319438 158080 319444 158092
rect 286928 158052 319444 158080
rect 286928 158040 286934 158052
rect 319438 158040 319444 158052
rect 319496 158040 319502 158092
rect 398466 158040 398472 158092
rect 398524 158080 398530 158092
rect 441706 158080 441712 158092
rect 398524 158052 441712 158080
rect 398524 158040 398530 158052
rect 441706 158040 441712 158052
rect 441764 158040 441770 158092
rect 275830 157972 275836 158024
rect 275888 158012 275894 158024
rect 333606 158012 333612 158024
rect 275888 157984 333612 158012
rect 275888 157972 275894 157984
rect 333606 157972 333612 157984
rect 333664 157972 333670 158024
rect 401042 157972 401048 158024
rect 401100 158012 401106 158024
rect 441798 158012 441804 158024
rect 401100 157984 441804 158012
rect 401100 157972 401106 157984
rect 441798 157972 441804 157984
rect 441856 157972 441862 158024
rect 159634 157904 159640 157956
rect 159692 157944 159698 157956
rect 285122 157944 285128 157956
rect 159692 157916 285128 157944
rect 159692 157904 159698 157916
rect 285122 157904 285128 157916
rect 285180 157904 285186 157956
rect 288250 157904 288256 157956
rect 288308 157944 288314 157956
rect 320542 157944 320548 157956
rect 288308 157916 320548 157944
rect 288308 157904 288314 157916
rect 320542 157904 320548 157916
rect 320600 157904 320606 157956
rect 403986 157904 403992 157956
rect 404044 157944 404050 157956
rect 438210 157944 438216 157956
rect 404044 157916 438216 157944
rect 404044 157904 404050 157916
rect 438210 157904 438216 157916
rect 438268 157904 438274 157956
rect 188706 157836 188712 157888
rect 188764 157876 188770 157888
rect 238478 157876 238484 157888
rect 188764 157848 238484 157876
rect 188764 157836 188770 157848
rect 238478 157836 238484 157848
rect 238536 157836 238542 157888
rect 290734 157836 290740 157888
rect 290792 157876 290798 157888
rect 321646 157876 321652 157888
rect 290792 157848 321652 157876
rect 290792 157836 290798 157848
rect 321646 157836 321652 157848
rect 321704 157836 321710 157888
rect 406470 157836 406476 157888
rect 406528 157876 406534 157888
rect 439682 157876 439688 157888
rect 406528 157848 439688 157876
rect 406528 157836 406534 157848
rect 439682 157836 439688 157848
rect 439740 157836 439746 157888
rect 206002 157768 206008 157820
rect 206060 157808 206066 157820
rect 238386 157808 238392 157820
rect 206060 157780 238392 157808
rect 206060 157768 206066 157780
rect 238386 157768 238392 157780
rect 238444 157768 238450 157820
rect 119890 157700 119896 157752
rect 119948 157740 119954 157752
rect 286134 157740 286140 157752
rect 119948 157712 286140 157740
rect 119948 157700 119954 157712
rect 286134 157700 286140 157712
rect 286192 157700 286198 157752
rect 97718 157632 97724 157684
rect 97776 157672 97782 157684
rect 297450 157672 297456 157684
rect 97776 157644 297456 157672
rect 97776 157632 97782 157644
rect 297450 157632 297456 157644
rect 297508 157632 297514 157684
rect 130562 157564 130568 157616
rect 130620 157604 130626 157616
rect 299382 157604 299388 157616
rect 130620 157576 299388 157604
rect 130620 157564 130626 157576
rect 299382 157564 299388 157576
rect 299440 157564 299446 157616
rect 331306 157496 331312 157548
rect 331364 157536 331370 157548
rect 354398 157536 354404 157548
rect 331364 157508 354404 157536
rect 331364 157496 331370 157508
rect 354398 157496 354404 157508
rect 354456 157496 354462 157548
rect 329742 157428 329748 157480
rect 329800 157468 329806 157480
rect 356974 157468 356980 157480
rect 329800 157440 356980 157468
rect 329800 157428 329806 157440
rect 356974 157428 356980 157440
rect 357032 157428 357038 157480
rect 327258 157360 327264 157412
rect 327316 157400 327322 157412
rect 355226 157400 355232 157412
rect 327316 157372 355232 157400
rect 327316 157360 327322 157372
rect 355226 157360 355232 157372
rect 355284 157360 355290 157412
rect 116210 157292 116216 157344
rect 116268 157332 116274 157344
rect 283742 157332 283748 157344
rect 116268 157304 283748 157332
rect 116268 157292 116274 157304
rect 283742 157292 283748 157304
rect 283800 157332 283806 157344
rect 284018 157332 284024 157344
rect 283800 157304 284024 157332
rect 283800 157292 283806 157304
rect 284018 157292 284024 157304
rect 284076 157292 284082 157344
rect 284478 157292 284484 157344
rect 284536 157332 284542 157344
rect 285582 157332 285588 157344
rect 284536 157304 285588 157332
rect 284536 157292 284542 157304
rect 285582 157292 285588 157304
rect 285640 157332 285646 157344
rect 347590 157332 347596 157344
rect 285640 157304 347596 157332
rect 285640 157292 285646 157304
rect 347590 157292 347596 157304
rect 347648 157292 347654 157344
rect 118234 157224 118240 157276
rect 118292 157264 118298 157276
rect 285398 157264 285404 157276
rect 118292 157236 285404 157264
rect 118292 157224 118298 157236
rect 285398 157224 285404 157236
rect 285456 157264 285462 157276
rect 290918 157264 290924 157276
rect 285456 157236 290924 157264
rect 285456 157224 285462 157236
rect 290918 157224 290924 157236
rect 290976 157224 290982 157276
rect 282546 157196 282552 157208
rect 277366 157168 282552 157196
rect 135898 156952 135904 157004
rect 135956 156992 135962 157004
rect 277366 156992 277394 157168
rect 282546 157156 282552 157168
rect 282604 157196 282610 157208
rect 335814 157196 335820 157208
rect 282604 157168 335820 157196
rect 282604 157156 282610 157168
rect 335814 157156 335820 157168
rect 335872 157156 335878 157208
rect 280062 157088 280068 157140
rect 280120 157128 280126 157140
rect 339310 157128 339316 157140
rect 280120 157100 339316 157128
rect 280120 157088 280126 157100
rect 339310 157088 339316 157100
rect 339368 157088 339374 157140
rect 278590 157020 278596 157072
rect 278648 157060 278654 157072
rect 330294 157060 330300 157072
rect 278648 157032 330300 157060
rect 278648 157020 278654 157032
rect 330294 157020 330300 157032
rect 330352 157020 330358 157072
rect 282822 156992 282828 157004
rect 135956 156964 277394 156992
rect 282380 156964 282828 156992
rect 135956 156952 135962 156964
rect 137002 156884 137008 156936
rect 137060 156924 137066 156936
rect 282380 156924 282408 156964
rect 282822 156952 282828 156964
rect 282880 156992 282886 157004
rect 336918 156992 336924 157004
rect 282880 156964 336924 156992
rect 282880 156952 282886 156964
rect 336918 156952 336924 156964
rect 336976 156952 336982 157004
rect 137060 156896 282408 156924
rect 137060 156884 137066 156896
rect 286134 156884 286140 156936
rect 286192 156924 286198 156936
rect 286962 156924 286968 156936
rect 286192 156896 286968 156924
rect 286192 156884 286198 156896
rect 286962 156884 286968 156896
rect 287020 156924 287026 156936
rect 334526 156924 334532 156936
rect 287020 156896 334532 156924
rect 287020 156884 287026 156896
rect 334526 156884 334532 156896
rect 334584 156884 334590 156936
rect 138382 156816 138388 156868
rect 138440 156856 138446 156868
rect 279970 156856 279976 156868
rect 138440 156828 279976 156856
rect 138440 156816 138446 156828
rect 279970 156816 279976 156828
rect 280028 156816 280034 156868
rect 283742 156816 283748 156868
rect 283800 156856 283806 156868
rect 316034 156856 316040 156868
rect 283800 156828 316040 156856
rect 283800 156816 283806 156828
rect 316034 156816 316040 156828
rect 316092 156816 316098 156868
rect 139670 156748 139676 156800
rect 139728 156788 139734 156800
rect 280062 156788 280068 156800
rect 139728 156760 280068 156788
rect 139728 156748 139734 156760
rect 280062 156748 280068 156760
rect 280120 156748 280126 156800
rect 290642 156748 290648 156800
rect 290700 156788 290706 156800
rect 323118 156788 323124 156800
rect 290700 156760 323124 156788
rect 290700 156748 290706 156760
rect 323118 156748 323124 156760
rect 323176 156748 323182 156800
rect 282914 156680 282920 156732
rect 282972 156720 282978 156732
rect 284110 156720 284116 156732
rect 282972 156692 284116 156720
rect 282972 156680 282978 156692
rect 284110 156680 284116 156692
rect 284168 156720 284174 156732
rect 317046 156720 317052 156732
rect 284168 156692 317052 156720
rect 284168 156680 284174 156692
rect 317046 156680 317052 156692
rect 317104 156680 317110 156732
rect 125594 156612 125600 156664
rect 125652 156652 125658 156664
rect 252830 156652 252836 156664
rect 125652 156624 252836 156652
rect 125652 156612 125658 156624
rect 252830 156612 252836 156624
rect 252888 156612 252894 156664
rect 253290 156612 253296 156664
rect 253348 156652 253354 156664
rect 275002 156652 275008 156664
rect 253348 156624 275008 156652
rect 253348 156612 253354 156624
rect 275002 156612 275008 156624
rect 275060 156612 275066 156664
rect 290182 156612 290188 156664
rect 290240 156652 290246 156664
rect 331214 156652 331220 156664
rect 290240 156624 331220 156652
rect 290240 156612 290246 156624
rect 331214 156612 331220 156624
rect 331272 156612 331278 156664
rect 184014 156544 184020 156596
rect 184072 156584 184078 156596
rect 280982 156584 280988 156596
rect 184072 156556 280988 156584
rect 184072 156544 184078 156556
rect 280982 156544 280988 156556
rect 281040 156544 281046 156596
rect 287514 156544 287520 156596
rect 287572 156584 287578 156596
rect 313274 156584 313280 156596
rect 287572 156556 313280 156584
rect 287572 156544 287578 156556
rect 313274 156544 313280 156556
rect 313332 156544 313338 156596
rect 185946 156476 185952 156528
rect 186004 156516 186010 156528
rect 280890 156516 280896 156528
rect 186004 156488 280896 156516
rect 186004 156476 186010 156488
rect 280890 156476 280896 156488
rect 280948 156476 280954 156528
rect 285950 156476 285956 156528
rect 286008 156516 286014 156528
rect 302234 156516 302240 156528
rect 286008 156488 302240 156516
rect 286008 156476 286014 156488
rect 302234 156476 302240 156488
rect 302292 156476 302298 156528
rect 191466 156408 191472 156460
rect 191524 156448 191530 156460
rect 280798 156448 280804 156460
rect 191524 156420 280804 156448
rect 191524 156408 191530 156420
rect 280798 156408 280804 156420
rect 280856 156408 280862 156460
rect 279970 156340 279976 156392
rect 280028 156380 280034 156392
rect 338114 156380 338120 156392
rect 280028 156352 338120 156380
rect 280028 156340 280034 156352
rect 338114 156340 338120 156352
rect 338172 156340 338178 156392
rect 123938 156272 123944 156324
rect 123996 156312 124002 156324
rect 290642 156312 290648 156324
rect 123996 156284 290648 156312
rect 123996 156272 124002 156284
rect 290642 156272 290648 156284
rect 290700 156272 290706 156324
rect 134610 156204 134616 156256
rect 134668 156244 134674 156256
rect 286134 156244 286140 156256
rect 134668 156216 286140 156244
rect 134668 156204 134674 156216
rect 286134 156204 286140 156216
rect 286192 156204 286198 156256
rect 117314 156136 117320 156188
rect 117372 156176 117378 156188
rect 282914 156176 282920 156188
rect 117372 156148 282920 156176
rect 117372 156136 117378 156148
rect 282914 156136 282920 156148
rect 282972 156136 282978 156188
rect 148686 156068 148692 156120
rect 148744 156108 148750 156120
rect 284478 156108 284484 156120
rect 148744 156080 284484 156108
rect 148744 156068 148750 156080
rect 284478 156068 284484 156080
rect 284536 156068 284542 156120
rect 271138 155864 271144 155916
rect 271196 155904 271202 155916
rect 276382 155904 276388 155916
rect 271196 155876 276388 155904
rect 271196 155864 271202 155876
rect 276382 155864 276388 155876
rect 276440 155864 276446 155916
rect 283558 155864 283564 155916
rect 283616 155904 283622 155916
rect 285950 155904 285956 155916
rect 283616 155876 285956 155904
rect 283616 155864 283622 155876
rect 285950 155864 285956 155876
rect 286008 155864 286014 155916
rect 286134 155864 286140 155916
rect 286192 155904 286198 155916
rect 345106 155904 345112 155916
rect 286192 155876 345112 155904
rect 286192 155864 286198 155876
rect 345106 155864 345112 155876
rect 345164 155864 345170 155916
rect 276014 155796 276020 155848
rect 276072 155836 276078 155848
rect 277210 155836 277216 155848
rect 276072 155808 277216 155836
rect 276072 155796 276078 155808
rect 277210 155796 277216 155808
rect 277268 155836 277274 155848
rect 346394 155836 346400 155848
rect 277268 155808 346400 155836
rect 277268 155796 277274 155808
rect 346394 155796 346400 155808
rect 346452 155796 346458 155848
rect 141786 155728 141792 155780
rect 141844 155768 141850 155780
rect 285490 155768 285496 155780
rect 141844 155740 285496 155768
rect 141844 155728 141850 155740
rect 285490 155728 285496 155740
rect 285548 155768 285554 155780
rect 341150 155768 341156 155780
rect 285548 155740 341156 155768
rect 285548 155728 285554 155740
rect 341150 155728 341156 155740
rect 341208 155728 341214 155780
rect 282362 155660 282368 155712
rect 282420 155700 282426 155712
rect 282638 155700 282644 155712
rect 282420 155672 282644 155700
rect 282420 155660 282426 155672
rect 282638 155660 282644 155672
rect 282696 155700 282702 155712
rect 348694 155700 348700 155712
rect 282696 155672 348700 155700
rect 282696 155660 282702 155672
rect 348694 155660 348700 155672
rect 348752 155660 348758 155712
rect 143074 155592 143080 155644
rect 143132 155632 143138 155644
rect 282730 155632 282736 155644
rect 143132 155604 282736 155632
rect 143132 155592 143138 155604
rect 282730 155592 282736 155604
rect 282788 155632 282794 155644
rect 342346 155632 342352 155644
rect 282788 155604 342352 155632
rect 282788 155592 282794 155604
rect 342346 155592 342352 155604
rect 342404 155592 342410 155644
rect 140682 155524 140688 155576
rect 140740 155564 140746 155576
rect 279602 155564 279608 155576
rect 140740 155536 279608 155564
rect 140740 155524 140746 155536
rect 279602 155524 279608 155536
rect 279660 155564 279666 155576
rect 339586 155564 339592 155576
rect 279660 155536 339592 155564
rect 279660 155524 279666 155536
rect 339586 155524 339592 155536
rect 339644 155524 339650 155576
rect 148778 155456 148784 155508
rect 148836 155496 148842 155508
rect 282362 155496 282368 155508
rect 148836 155468 282368 155496
rect 148836 155456 148842 155468
rect 282362 155456 282368 155468
rect 282420 155456 282426 155508
rect 282914 155456 282920 155508
rect 282972 155496 282978 155508
rect 284202 155496 284208 155508
rect 282972 155468 284208 155496
rect 282972 155456 282978 155468
rect 284202 155456 284208 155468
rect 284260 155496 284266 155508
rect 343910 155496 343916 155508
rect 284260 155468 343916 155496
rect 284260 155456 284266 155468
rect 343910 155456 343916 155468
rect 343968 155456 343974 155508
rect 145282 155388 145288 155440
rect 145340 155428 145346 155440
rect 279694 155428 279700 155440
rect 145340 155400 279700 155428
rect 145340 155388 145346 155400
rect 279694 155388 279700 155400
rect 279752 155428 279758 155440
rect 286134 155428 286140 155440
rect 279752 155400 286140 155428
rect 279752 155388 279758 155400
rect 286134 155388 286140 155400
rect 286192 155388 286198 155440
rect 289538 155388 289544 155440
rect 289596 155428 289602 155440
rect 324222 155428 324228 155440
rect 289596 155400 324228 155428
rect 289596 155388 289602 155400
rect 324222 155388 324228 155400
rect 324280 155388 324286 155440
rect 146386 155320 146392 155372
rect 146444 155360 146450 155372
rect 276014 155360 276020 155372
rect 146444 155332 276020 155360
rect 146444 155320 146450 155332
rect 276014 155320 276020 155332
rect 276072 155320 276078 155372
rect 299382 155320 299388 155372
rect 299440 155360 299446 155372
rect 327258 155360 327264 155372
rect 299440 155332 327264 155360
rect 299440 155320 299446 155332
rect 327258 155320 327264 155332
rect 327316 155320 327322 155372
rect 148410 155252 148416 155304
rect 148468 155292 148474 155304
rect 269942 155292 269948 155304
rect 148468 155264 269948 155292
rect 148468 155252 148474 155264
rect 269942 155252 269948 155264
rect 270000 155252 270006 155304
rect 288894 155252 288900 155304
rect 288952 155292 288958 155304
rect 320174 155292 320180 155304
rect 288952 155264 320180 155292
rect 288952 155252 288958 155264
rect 320174 155252 320180 155264
rect 320232 155252 320238 155304
rect 150986 155184 150992 155236
rect 151044 155224 151050 155236
rect 270034 155224 270040 155236
rect 151044 155196 270040 155224
rect 151044 155184 151050 155196
rect 270034 155184 270040 155196
rect 270092 155184 270098 155236
rect 291654 155184 291660 155236
rect 291712 155224 291718 155236
rect 338114 155224 338120 155236
rect 291712 155196 338120 155224
rect 291712 155184 291718 155196
rect 338114 155184 338120 155196
rect 338172 155184 338178 155236
rect 201034 155116 201040 155168
rect 201092 155156 201098 155168
rect 275370 155156 275376 155168
rect 201092 155128 275376 155156
rect 201092 155116 201098 155128
rect 275370 155116 275376 155128
rect 275428 155116 275434 155168
rect 286042 155116 286048 155168
rect 286100 155156 286106 155168
rect 306374 155156 306380 155168
rect 286100 155128 306380 155156
rect 286100 155116 286106 155128
rect 306374 155116 306380 155128
rect 306432 155116 306438 155168
rect 203426 155048 203432 155100
rect 203484 155088 203490 155100
rect 275462 155088 275468 155100
rect 203484 155060 275468 155088
rect 203484 155048 203490 155060
rect 275462 155048 275468 155060
rect 275520 155048 275526 155100
rect 229094 154980 229100 155032
rect 229152 155020 229158 155032
rect 272242 155020 272248 155032
rect 229152 154992 272248 155020
rect 229152 154980 229158 154992
rect 272242 154980 272248 154992
rect 272300 154980 272306 155032
rect 155770 154912 155776 154964
rect 155828 154952 155834 154964
rect 298370 154952 298376 154964
rect 155828 154924 298376 154952
rect 155828 154912 155834 154924
rect 298370 154912 298376 154924
rect 298428 154952 298434 154964
rect 299382 154952 299388 154964
rect 298428 154924 299388 154952
rect 298428 154912 298434 154924
rect 299382 154912 299388 154924
rect 299440 154912 299446 154964
rect 124766 154844 124772 154896
rect 124824 154884 124830 154896
rect 289538 154884 289544 154896
rect 124824 154856 289544 154884
rect 124824 154844 124830 154856
rect 289538 154844 289544 154856
rect 289596 154844 289602 154896
rect 143994 154776 144000 154828
rect 144052 154816 144058 154828
rect 282914 154816 282920 154828
rect 144052 154788 282920 154816
rect 144052 154776 144058 154788
rect 282914 154776 282920 154788
rect 282972 154776 282978 154828
rect 125410 154504 125416 154556
rect 125468 154544 125474 154556
rect 276014 154544 276020 154556
rect 125468 154516 276020 154544
rect 125468 154504 125474 154516
rect 276014 154504 276020 154516
rect 276072 154504 276078 154556
rect 279786 154504 279792 154556
rect 279844 154544 279850 154556
rect 280062 154544 280068 154556
rect 279844 154516 280068 154544
rect 279844 154504 279850 154516
rect 280062 154504 280068 154516
rect 280120 154544 280126 154556
rect 351086 154544 351092 154556
rect 280120 154516 351092 154544
rect 280120 154504 280126 154516
rect 351086 154504 351092 154516
rect 351144 154504 351150 154556
rect 153838 154436 153844 154488
rect 153896 154476 153902 154488
rect 297910 154476 297916 154488
rect 153896 154448 297916 154476
rect 153896 154436 153902 154448
rect 297910 154436 297916 154448
rect 297968 154476 297974 154488
rect 353294 154476 353300 154488
rect 297968 154448 353300 154476
rect 297968 154436 297974 154448
rect 353294 154436 353300 154448
rect 353352 154436 353358 154488
rect 152642 154368 152648 154420
rect 152700 154408 152706 154420
rect 152700 154380 277394 154408
rect 152700 154368 152706 154380
rect 141510 154300 141516 154352
rect 141568 154340 141574 154352
rect 272518 154340 272524 154352
rect 141568 154312 272524 154340
rect 141568 154300 141574 154312
rect 272518 154300 272524 154312
rect 272576 154300 272582 154352
rect 277366 154340 277394 154380
rect 290826 154368 290832 154420
rect 290884 154408 290890 154420
rect 345750 154408 345756 154420
rect 290884 154380 345756 154408
rect 290884 154368 290890 154380
rect 345750 154368 345756 154380
rect 345808 154368 345814 154420
rect 281350 154340 281356 154352
rect 277366 154312 281356 154340
rect 281350 154300 281356 154312
rect 281408 154340 281414 154352
rect 352190 154340 352196 154352
rect 281408 154312 352196 154340
rect 281408 154300 281414 154312
rect 352190 154300 352196 154312
rect 352248 154300 352254 154352
rect 149882 154232 149888 154284
rect 149940 154272 149946 154284
rect 279878 154272 279884 154284
rect 149940 154244 279884 154272
rect 149940 154232 149946 154244
rect 279878 154232 279884 154244
rect 279936 154272 279942 154284
rect 349798 154272 349804 154284
rect 279936 154244 349804 154272
rect 279936 154232 279942 154244
rect 349798 154232 349804 154244
rect 349856 154232 349862 154284
rect 276014 154164 276020 154216
rect 276072 154204 276078 154216
rect 277302 154204 277308 154216
rect 276072 154176 277308 154204
rect 276072 154164 276078 154176
rect 277302 154164 277308 154176
rect 277360 154204 277366 154216
rect 324866 154204 324872 154216
rect 277360 154176 324872 154204
rect 277360 154164 277366 154176
rect 324866 154164 324872 154176
rect 324924 154164 324930 154216
rect 151354 154096 151360 154148
rect 151412 154136 151418 154148
rect 280062 154136 280068 154148
rect 151412 154108 280068 154136
rect 151412 154096 151418 154108
rect 280062 154096 280068 154108
rect 280120 154096 280126 154148
rect 329742 154136 329748 154148
rect 287026 154108 329748 154136
rect 157058 154028 157064 154080
rect 157116 154068 157122 154080
rect 283926 154068 283932 154080
rect 157116 154040 283932 154068
rect 157116 154028 157122 154040
rect 283926 154028 283932 154040
rect 283984 154068 283990 154080
rect 287026 154068 287054 154108
rect 329742 154096 329748 154108
rect 329800 154096 329806 154148
rect 283984 154040 287054 154068
rect 283984 154028 283990 154040
rect 297450 154028 297456 154080
rect 297508 154068 297514 154080
rect 331306 154068 331312 154080
rect 297508 154040 331312 154068
rect 297508 154028 297514 154040
rect 331306 154028 331312 154040
rect 331364 154028 331370 154080
rect 146018 153960 146024 154012
rect 146076 154000 146082 154012
rect 269850 154000 269856 154012
rect 146076 153972 269856 154000
rect 146076 153960 146082 153972
rect 269850 153960 269856 153972
rect 269908 153960 269914 154012
rect 195882 153892 195888 153944
rect 195940 153932 195946 153944
rect 278130 153932 278136 153944
rect 195940 153904 278136 153932
rect 195940 153892 195946 153904
rect 278130 153892 278136 153904
rect 278188 153892 278194 153944
rect 164234 153824 164240 153876
rect 164292 153864 164298 153876
rect 259914 153864 259920 153876
rect 164292 153836 259920 153864
rect 164292 153824 164298 153836
rect 259914 153824 259920 153836
rect 259972 153824 259978 153876
rect 287422 153824 287428 153876
rect 287480 153864 287486 153876
rect 316034 153864 316040 153876
rect 287480 153836 316040 153864
rect 287480 153824 287486 153836
rect 316034 153824 316040 153836
rect 316092 153824 316098 153876
rect 198458 153756 198464 153808
rect 198516 153796 198522 153808
rect 278222 153796 278228 153808
rect 198516 153768 278228 153796
rect 198516 153756 198522 153768
rect 278222 153756 278228 153768
rect 278280 153756 278286 153808
rect 202874 153688 202880 153740
rect 202932 153728 202938 153740
rect 266814 153728 266820 153740
rect 202932 153700 266820 153728
rect 202932 153688 202938 153700
rect 266814 153688 266820 153700
rect 266872 153688 266878 153740
rect 231854 153620 231860 153672
rect 231912 153660 231918 153672
rect 272150 153660 272156 153672
rect 231912 153632 272156 153660
rect 231912 153620 231918 153632
rect 272150 153620 272156 153632
rect 272208 153620 272214 153672
rect 154482 153552 154488 153604
rect 154540 153592 154546 153604
rect 296714 153592 296720 153604
rect 154540 153564 296720 153592
rect 154540 153552 154546 153564
rect 296714 153552 296720 153564
rect 296772 153592 296778 153604
rect 297450 153592 297456 153604
rect 296772 153564 297456 153592
rect 296772 153552 296778 153564
rect 297450 153552 297456 153564
rect 297508 153552 297514 153604
rect 233234 152668 233240 152720
rect 233292 152708 233298 152720
rect 272058 152708 272064 152720
rect 233292 152680 272064 152708
rect 233292 152668 233298 152680
rect 272058 152668 272064 152680
rect 272116 152668 272122 152720
rect 227714 152600 227720 152652
rect 227772 152640 227778 152652
rect 269758 152640 269764 152652
rect 227772 152612 269764 152640
rect 227772 152600 227778 152612
rect 269758 152600 269764 152612
rect 269816 152600 269822 152652
rect 288802 152600 288808 152652
rect 288860 152640 288866 152652
rect 324314 152640 324320 152652
rect 288860 152612 324320 152640
rect 288860 152600 288866 152612
rect 324314 152600 324320 152612
rect 324372 152600 324378 152652
rect 193214 152532 193220 152584
rect 193272 152572 193278 152584
rect 265434 152572 265440 152584
rect 193272 152544 265440 152572
rect 193272 152532 193278 152544
rect 265434 152532 265440 152544
rect 265492 152532 265498 152584
rect 294322 152532 294328 152584
rect 294380 152572 294386 152584
rect 349154 152572 349160 152584
rect 294380 152544 349160 152572
rect 294380 152532 294386 152544
rect 349154 152532 349160 152544
rect 349212 152532 349218 152584
rect 168374 152464 168380 152516
rect 168432 152504 168438 152516
rect 242250 152504 242256 152516
rect 168432 152476 242256 152504
rect 168432 152464 168438 152476
rect 242250 152464 242256 152476
rect 242308 152464 242314 152516
rect 299106 152464 299112 152516
rect 299164 152504 299170 152516
rect 376754 152504 376760 152516
rect 299164 152476 376760 152504
rect 299164 152464 299170 152476
rect 376754 152464 376760 152476
rect 376812 152464 376818 152516
rect 272518 151784 272524 151836
rect 272576 151824 272582 151836
rect 278958 151824 278964 151836
rect 272576 151796 278964 151824
rect 272576 151784 272582 151796
rect 278958 151784 278964 151796
rect 279016 151784 279022 151836
rect 209774 151172 209780 151224
rect 209832 151212 209838 151224
rect 268102 151212 268108 151224
rect 209832 151184 268108 151212
rect 209832 151172 209838 151184
rect 268102 151172 268108 151184
rect 268160 151172 268166 151224
rect 284386 151172 284392 151224
rect 284444 151212 284450 151224
rect 299566 151212 299572 151224
rect 284444 151184 299572 151212
rect 284444 151172 284450 151184
rect 299566 151172 299572 151184
rect 299624 151172 299630 151224
rect 175274 151104 175280 151156
rect 175332 151144 175338 151156
rect 261478 151144 261484 151156
rect 175332 151116 261484 151144
rect 175332 151104 175338 151116
rect 261478 151104 261484 151116
rect 261536 151104 261542 151156
rect 290090 151104 290096 151156
rect 290148 151144 290154 151156
rect 324406 151144 324412 151156
rect 290148 151116 324412 151144
rect 290148 151104 290154 151116
rect 324406 151104 324412 151116
rect 324464 151104 324470 151156
rect 146294 151036 146300 151088
rect 146352 151076 146358 151088
rect 257154 151076 257160 151088
rect 146352 151048 257160 151076
rect 146352 151036 146358 151048
rect 257154 151036 257160 151048
rect 257212 151036 257218 151088
rect 292942 151036 292948 151088
rect 293000 151076 293006 151088
rect 340874 151076 340880 151088
rect 293000 151048 340880 151076
rect 293000 151036 293006 151048
rect 340874 151036 340880 151048
rect 340932 151036 340938 151088
rect 268194 150424 268200 150476
rect 268252 150464 268258 150476
rect 273898 150464 273904 150476
rect 268252 150436 273904 150464
rect 268252 150424 268258 150436
rect 273898 150424 273904 150436
rect 273956 150424 273962 150476
rect 213914 149812 213920 149864
rect 213972 149852 213978 149864
rect 269574 149852 269580 149864
rect 213972 149824 269580 149852
rect 213972 149812 213978 149824
rect 269574 149812 269580 149824
rect 269632 149812 269638 149864
rect 285858 149812 285864 149864
rect 285916 149852 285922 149864
rect 303614 149852 303620 149864
rect 285916 149824 303620 149852
rect 285916 149812 285922 149824
rect 303614 149812 303620 149824
rect 303672 149812 303678 149864
rect 184934 149744 184940 149796
rect 184992 149784 184998 149796
rect 264054 149784 264060 149796
rect 184992 149756 264060 149784
rect 184992 149744 184998 149756
rect 264054 149744 264060 149756
rect 264112 149744 264118 149796
rect 292850 149744 292856 149796
rect 292908 149784 292914 149796
rect 345014 149784 345020 149796
rect 292908 149756 345020 149784
rect 292908 149744 292914 149756
rect 345014 149744 345020 149756
rect 345072 149744 345078 149796
rect 157334 149676 157340 149728
rect 157392 149716 157398 149728
rect 258350 149716 258356 149728
rect 157392 149688 258356 149716
rect 157392 149676 157398 149688
rect 258350 149676 258356 149688
rect 258408 149676 258414 149728
rect 295702 149676 295708 149728
rect 295760 149716 295766 149728
rect 357434 149716 357440 149728
rect 295760 149688 357440 149716
rect 295760 149676 295766 149688
rect 357434 149676 357440 149688
rect 357492 149676 357498 149728
rect 215294 148452 215300 148504
rect 215352 148492 215358 148504
rect 269482 148492 269488 148504
rect 215352 148464 269488 148492
rect 215352 148452 215358 148464
rect 269482 148452 269488 148464
rect 269540 148452 269546 148504
rect 189074 148384 189080 148436
rect 189132 148424 189138 148436
rect 263962 148424 263968 148436
rect 189132 148396 263968 148424
rect 189132 148384 189138 148396
rect 263962 148384 263968 148396
rect 264020 148384 264026 148436
rect 291562 148384 291568 148436
rect 291620 148424 291626 148436
rect 332594 148424 332600 148436
rect 291620 148396 332600 148424
rect 291620 148384 291626 148396
rect 332594 148384 332600 148396
rect 332652 148384 332658 148436
rect 135254 148316 135260 148368
rect 135312 148356 135318 148368
rect 254210 148356 254216 148368
rect 135312 148328 254216 148356
rect 135312 148316 135318 148328
rect 254210 148316 254216 148328
rect 254268 148316 254274 148368
rect 294230 148316 294236 148368
rect 294288 148356 294294 148368
rect 351914 148356 351920 148368
rect 294288 148328 351920 148356
rect 294288 148316 294294 148328
rect 351914 148316 351920 148328
rect 351972 148316 351978 148368
rect 176654 146956 176660 147008
rect 176712 146996 176718 147008
rect 262490 146996 262496 147008
rect 176712 146968 262496 146996
rect 176712 146956 176718 146968
rect 262490 146956 262496 146968
rect 262548 146956 262554 147008
rect 287330 146956 287336 147008
rect 287388 146996 287394 147008
rect 310514 146996 310520 147008
rect 287388 146968 310520 146996
rect 287388 146956 287394 146968
rect 310514 146956 310520 146968
rect 310572 146956 310578 147008
rect 128354 146888 128360 146940
rect 128412 146928 128418 146940
rect 252738 146928 252744 146940
rect 128412 146900 252744 146928
rect 128412 146888 128418 146900
rect 252738 146888 252744 146900
rect 252796 146888 252802 146940
rect 253382 146888 253388 146940
rect 253440 146928 253446 146940
rect 273622 146928 273628 146940
rect 253440 146900 273628 146928
rect 253440 146888 253446 146900
rect 273622 146888 273628 146900
rect 273680 146888 273686 146940
rect 289998 146888 290004 146940
rect 290056 146928 290062 146940
rect 328454 146928 328460 146940
rect 290056 146900 328460 146928
rect 290056 146888 290062 146900
rect 328454 146888 328460 146900
rect 328512 146888 328518 146940
rect 279510 146548 279516 146600
rect 279568 146588 279574 146600
rect 280430 146588 280436 146600
rect 279568 146560 280436 146588
rect 279568 146548 279574 146560
rect 280430 146548 280436 146560
rect 280488 146548 280494 146600
rect 219434 145664 219440 145716
rect 219492 145704 219498 145716
rect 270862 145704 270868 145716
rect 219492 145676 270868 145704
rect 219492 145664 219498 145676
rect 270862 145664 270868 145676
rect 270920 145664 270926 145716
rect 287238 145664 287244 145716
rect 287296 145704 287302 145716
rect 314654 145704 314660 145716
rect 287296 145676 314660 145704
rect 287296 145664 287302 145676
rect 314654 145664 314660 145676
rect 314712 145664 314718 145716
rect 195974 145596 195980 145648
rect 196032 145636 196038 145648
rect 265342 145636 265348 145648
rect 196032 145608 265348 145636
rect 196032 145596 196038 145608
rect 265342 145596 265348 145608
rect 265400 145596 265406 145648
rect 292758 145596 292764 145648
rect 292816 145636 292822 145648
rect 342254 145636 342260 145648
rect 292816 145608 342260 145636
rect 292816 145596 292822 145608
rect 342254 145596 342260 145608
rect 342312 145596 342318 145648
rect 153194 145528 153200 145580
rect 153252 145568 153258 145580
rect 255958 145568 255964 145580
rect 153252 145540 255964 145568
rect 153252 145528 153258 145540
rect 255958 145528 255964 145540
rect 256016 145528 256022 145580
rect 265618 145528 265624 145580
rect 265676 145568 265682 145580
rect 274910 145568 274916 145580
rect 265676 145540 274916 145568
rect 265676 145528 265682 145540
rect 274910 145528 274916 145540
rect 274968 145528 274974 145580
rect 275002 145528 275008 145580
rect 275060 145568 275066 145580
rect 280338 145568 280344 145580
rect 275060 145540 280344 145568
rect 275060 145528 275066 145540
rect 280338 145528 280344 145540
rect 280396 145528 280402 145580
rect 283190 145528 283196 145580
rect 283248 145568 283254 145580
rect 287238 145568 287244 145580
rect 283248 145540 287244 145568
rect 283248 145528 283254 145540
rect 287238 145528 287244 145540
rect 287296 145528 287302 145580
rect 294138 145528 294144 145580
rect 294196 145568 294202 145580
rect 350534 145568 350540 145580
rect 294196 145540 350540 145568
rect 294196 145528 294202 145540
rect 350534 145528 350540 145540
rect 350592 145528 350598 145580
rect 218054 144304 218060 144356
rect 218112 144344 218118 144356
rect 269390 144344 269396 144356
rect 218112 144316 269396 144344
rect 218112 144304 218118 144316
rect 269390 144304 269396 144316
rect 269448 144304 269454 144356
rect 154574 144236 154580 144288
rect 154632 144276 154638 144288
rect 258258 144276 258264 144288
rect 154632 144248 258264 144276
rect 154632 144236 154638 144248
rect 258258 144236 258264 144248
rect 258316 144236 258322 144288
rect 288710 144236 288716 144288
rect 288768 144276 288774 144288
rect 317414 144276 317420 144288
rect 288768 144248 317420 144276
rect 288768 144236 288774 144248
rect 317414 144236 317420 144248
rect 317472 144236 317478 144288
rect 143534 144168 143540 144220
rect 143592 144208 143598 144220
rect 255774 144208 255780 144220
rect 143592 144180 255780 144208
rect 143592 144168 143598 144180
rect 255774 144168 255780 144180
rect 255832 144168 255838 144220
rect 294046 144168 294052 144220
rect 294104 144208 294110 144220
rect 353294 144208 353300 144220
rect 294104 144180 353300 144208
rect 294104 144168 294110 144180
rect 353294 144168 353300 144180
rect 353352 144168 353358 144220
rect 269758 144032 269764 144084
rect 269816 144072 269822 144084
rect 276290 144072 276296 144084
rect 269816 144044 276296 144072
rect 269816 144032 269822 144044
rect 276290 144032 276296 144044
rect 276348 144032 276354 144084
rect 235994 142944 236000 142996
rect 236052 142984 236058 142996
rect 273530 142984 273536 142996
rect 236052 142956 273536 142984
rect 236052 142944 236058 142956
rect 273530 142944 273536 142956
rect 273588 142944 273594 142996
rect 183554 142876 183560 142928
rect 183612 142916 183618 142928
rect 263870 142916 263876 142928
rect 183612 142888 263876 142916
rect 183612 142876 183618 142888
rect 263870 142876 263876 142888
rect 263928 142876 263934 142928
rect 288618 142876 288624 142928
rect 288676 142916 288682 142928
rect 321554 142916 321560 142928
rect 288676 142888 321560 142916
rect 288676 142876 288682 142888
rect 321554 142876 321560 142888
rect 321612 142876 321618 142928
rect 132494 142808 132500 142860
rect 132552 142848 132558 142860
rect 253198 142848 253204 142860
rect 132552 142820 253204 142848
rect 132552 142808 132558 142820
rect 253198 142808 253204 142820
rect 253256 142808 253262 142860
rect 295610 142808 295616 142860
rect 295668 142848 295674 142860
rect 360194 142848 360200 142860
rect 295668 142820 360200 142848
rect 295668 142808 295674 142820
rect 360194 142808 360200 142820
rect 360252 142808 360258 142860
rect 193306 141516 193312 141568
rect 193364 141556 193370 141568
rect 265250 141556 265256 141568
rect 193364 141528 265256 141556
rect 193364 141516 193370 141528
rect 265250 141516 265256 141528
rect 265308 141516 265314 141568
rect 139394 141448 139400 141500
rect 139452 141488 139458 141500
rect 254578 141488 254584 141500
rect 139452 141460 254584 141488
rect 139452 141448 139458 141460
rect 254578 141448 254584 141460
rect 254636 141448 254642 141500
rect 285766 141448 285772 141500
rect 285824 141488 285830 141500
rect 304994 141488 305000 141500
rect 285824 141460 305000 141488
rect 285824 141448 285830 141460
rect 304994 141448 305000 141460
rect 305052 141448 305058 141500
rect 121454 141380 121460 141432
rect 121512 141420 121518 141432
rect 251542 141420 251548 141432
rect 121512 141392 251548 141420
rect 121512 141380 121518 141392
rect 251542 141380 251548 141392
rect 251600 141380 251606 141432
rect 291470 141380 291476 141432
rect 291528 141420 291534 141432
rect 335354 141420 335360 141432
rect 291528 141392 335360 141420
rect 291528 141380 291534 141392
rect 335354 141380 335360 141392
rect 335412 141380 335418 141432
rect 197354 140156 197360 140208
rect 197412 140196 197418 140208
rect 266722 140196 266728 140208
rect 197412 140168 266728 140196
rect 197412 140156 197418 140168
rect 266722 140156 266728 140168
rect 266780 140156 266786 140208
rect 285030 140156 285036 140208
rect 285088 140196 285094 140208
rect 291470 140196 291476 140208
rect 285088 140168 291476 140196
rect 285088 140156 285094 140168
rect 291470 140156 291476 140168
rect 291528 140156 291534 140208
rect 150434 140088 150440 140140
rect 150492 140128 150498 140140
rect 257062 140128 257068 140140
rect 150492 140100 257068 140128
rect 150492 140088 150498 140100
rect 257062 140088 257068 140100
rect 257120 140088 257126 140140
rect 114554 140020 114560 140072
rect 114612 140060 114618 140072
rect 243630 140060 243636 140072
rect 114612 140032 243636 140060
rect 114612 140020 114618 140032
rect 243630 140020 243636 140032
rect 243688 140020 243694 140072
rect 291378 140020 291384 140072
rect 291436 140060 291442 140072
rect 339494 140060 339500 140072
rect 291436 140032 339500 140060
rect 291436 140020 291442 140032
rect 339494 140020 339500 140032
rect 339552 140020 339558 140072
rect 201494 138728 201500 138780
rect 201552 138768 201558 138780
rect 266630 138768 266636 138780
rect 201552 138740 266636 138768
rect 201552 138728 201558 138740
rect 266630 138728 266636 138740
rect 266688 138728 266694 138780
rect 126974 138660 126980 138712
rect 127032 138700 127038 138712
rect 252646 138700 252652 138712
rect 127032 138672 252652 138700
rect 127032 138660 127038 138672
rect 252646 138660 252652 138672
rect 252704 138660 252710 138712
rect 292666 138660 292672 138712
rect 292724 138700 292730 138712
rect 346394 138700 346400 138712
rect 292724 138672 346400 138700
rect 292724 138660 292730 138672
rect 346394 138660 346400 138672
rect 346452 138660 346458 138712
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 80698 137952 80704 137964
rect 3568 137924 80704 137952
rect 3568 137912 3574 137924
rect 80698 137912 80704 137924
rect 80756 137912 80762 137964
rect 211154 137368 211160 137420
rect 211212 137408 211218 137420
rect 268010 137408 268016 137420
rect 211212 137380 268016 137408
rect 211212 137368 211218 137380
rect 268010 137368 268016 137380
rect 268068 137368 268074 137420
rect 161474 137300 161480 137352
rect 161532 137340 161538 137352
rect 259822 137340 259828 137352
rect 161532 137312 259828 137340
rect 161532 137300 161538 137312
rect 259822 137300 259828 137312
rect 259880 137300 259886 137352
rect 107654 137232 107660 137284
rect 107712 137272 107718 137284
rect 246482 137272 246488 137284
rect 107712 137244 246488 137272
rect 107712 137232 107718 137244
rect 246482 137232 246488 137244
rect 246540 137232 246546 137284
rect 293954 137232 293960 137284
rect 294012 137272 294018 137284
rect 349246 137272 349252 137284
rect 294012 137244 349252 137272
rect 294012 137232 294018 137244
rect 349246 137232 349252 137244
rect 349304 137232 349310 137284
rect 222194 136008 222200 136060
rect 222252 136048 222258 136060
rect 270770 136048 270776 136060
rect 222252 136020 270776 136048
rect 222252 136008 222258 136020
rect 270770 136008 270776 136020
rect 270828 136008 270834 136060
rect 165614 135940 165620 135992
rect 165672 135980 165678 135992
rect 259730 135980 259736 135992
rect 165672 135952 259736 135980
rect 165672 135940 165678 135952
rect 259730 135940 259736 135952
rect 259788 135940 259794 135992
rect 103514 135872 103520 135924
rect 103572 135912 103578 135924
rect 248690 135912 248696 135924
rect 103572 135884 248696 135912
rect 103572 135872 103578 135884
rect 248690 135872 248696 135884
rect 248748 135872 248754 135924
rect 168466 134580 168472 134632
rect 168524 134620 168530 134632
rect 261294 134620 261300 134632
rect 168524 134592 261300 134620
rect 168524 134580 168530 134592
rect 261294 134580 261300 134592
rect 261352 134580 261358 134632
rect 147674 134512 147680 134564
rect 147732 134552 147738 134564
rect 256970 134552 256976 134564
rect 147732 134524 256976 134552
rect 147732 134512 147738 134524
rect 256970 134512 256976 134524
rect 257028 134512 257034 134564
rect 288526 134512 288532 134564
rect 288584 134552 288590 134564
rect 318794 134552 318800 134564
rect 288584 134524 318800 134552
rect 288584 134512 288590 134524
rect 318794 134512 318800 134524
rect 318852 134512 318858 134564
rect 191834 133220 191840 133272
rect 191892 133260 191898 133272
rect 265158 133260 265164 133272
rect 191892 133232 265164 133260
rect 191892 133220 191898 133232
rect 265158 133220 265164 133232
rect 265216 133220 265222 133272
rect 172514 133152 172520 133204
rect 172572 133192 172578 133204
rect 261202 133192 261208 133204
rect 172572 133164 261208 133192
rect 172572 133152 172578 133164
rect 261202 133152 261208 133164
rect 261260 133152 261266 133204
rect 261478 133152 261484 133204
rect 261536 133192 261542 133204
rect 276198 133192 276204 133204
rect 261536 133164 276204 133192
rect 261536 133152 261542 133164
rect 276198 133152 276204 133164
rect 276256 133152 276262 133204
rect 216674 131860 216680 131912
rect 216732 131900 216738 131912
rect 269298 131900 269304 131912
rect 216732 131872 269304 131900
rect 216732 131860 216738 131872
rect 269298 131860 269304 131872
rect 269356 131860 269362 131912
rect 179414 131792 179420 131844
rect 179472 131832 179478 131844
rect 262398 131832 262404 131844
rect 179472 131804 262404 131832
rect 179472 131792 179478 131804
rect 262398 131792 262404 131804
rect 262456 131792 262462 131844
rect 110414 131724 110420 131776
rect 110472 131764 110478 131776
rect 249978 131764 249984 131776
rect 110472 131736 249984 131764
rect 110472 131724 110478 131736
rect 249978 131724 249984 131736
rect 250036 131724 250042 131776
rect 288434 131724 288440 131776
rect 288492 131764 288498 131776
rect 322934 131764 322940 131776
rect 288492 131736 322940 131764
rect 288492 131724 288498 131736
rect 322934 131724 322940 131736
rect 322992 131724 322998 131776
rect 230474 130500 230480 130552
rect 230532 130540 230538 130552
rect 271966 130540 271972 130552
rect 230532 130512 271972 130540
rect 230532 130500 230538 130512
rect 271966 130500 271972 130512
rect 272024 130500 272030 130552
rect 186314 130432 186320 130484
rect 186372 130472 186378 130484
rect 263778 130472 263784 130484
rect 186372 130444 263784 130472
rect 186372 130432 186378 130444
rect 263778 130432 263784 130444
rect 263836 130432 263842 130484
rect 100754 130364 100760 130416
rect 100812 130404 100818 130416
rect 247770 130404 247776 130416
rect 100812 130376 247776 130404
rect 100812 130364 100818 130376
rect 247770 130364 247776 130376
rect 247828 130364 247834 130416
rect 289906 130364 289912 130416
rect 289964 130404 289970 130416
rect 325694 130404 325700 130416
rect 289964 130376 325700 130404
rect 289964 130364 289970 130376
rect 325694 130364 325700 130376
rect 325752 130364 325758 130416
rect 190454 129072 190460 129124
rect 190512 129112 190518 129124
rect 265066 129112 265072 129124
rect 190512 129084 265072 129112
rect 190512 129072 190518 129084
rect 265066 129072 265072 129084
rect 265124 129072 265130 129124
rect 149054 129004 149060 129056
rect 149112 129044 149118 129056
rect 256878 129044 256884 129056
rect 149112 129016 256884 129044
rect 149112 129004 149118 129016
rect 256878 129004 256884 129016
rect 256936 129004 256942 129056
rect 291286 129004 291292 129056
rect 291344 129044 291350 129056
rect 332686 129044 332692 129056
rect 291344 129016 332692 129044
rect 291344 129004 291350 129016
rect 332686 129004 332692 129016
rect 332744 129004 332750 129056
rect 204254 127644 204260 127696
rect 204312 127684 204318 127696
rect 266538 127684 266544 127696
rect 204312 127656 266544 127684
rect 204312 127644 204318 127656
rect 266538 127644 266544 127656
rect 266596 127644 266602 127696
rect 131114 127576 131120 127628
rect 131172 127616 131178 127628
rect 254118 127616 254124 127628
rect 131172 127588 254124 127616
rect 131172 127576 131178 127588
rect 254118 127576 254124 127588
rect 254176 127576 254182 127628
rect 291194 127576 291200 127628
rect 291252 127616 291258 127628
rect 336734 127616 336740 127628
rect 291252 127588 336740 127616
rect 291252 127576 291258 127588
rect 336734 127576 336740 127588
rect 336792 127576 336798 127628
rect 208394 126284 208400 126336
rect 208452 126324 208458 126336
rect 267918 126324 267924 126336
rect 208452 126296 267924 126324
rect 208452 126284 208458 126296
rect 267918 126284 267924 126296
rect 267976 126284 267982 126336
rect 138014 126216 138020 126268
rect 138072 126256 138078 126268
rect 255682 126256 255688 126268
rect 138072 126228 255688 126256
rect 138072 126216 138078 126228
rect 255682 126216 255688 126228
rect 255740 126216 255746 126268
rect 294598 126216 294604 126268
rect 294656 126256 294662 126268
rect 340966 126256 340972 126268
rect 294656 126228 340972 126256
rect 294656 126216 294662 126228
rect 340966 126216 340972 126228
rect 341024 126216 341030 126268
rect 280338 125536 280344 125588
rect 280396 125576 280402 125588
rect 281902 125576 281908 125588
rect 280396 125548 281908 125576
rect 280396 125536 280402 125548
rect 281902 125536 281908 125548
rect 281960 125536 281966 125588
rect 218146 124924 218152 124976
rect 218204 124964 218210 124976
rect 269206 124964 269212 124976
rect 218204 124936 269212 124964
rect 218204 124924 218210 124936
rect 269206 124924 269212 124936
rect 269264 124924 269270 124976
rect 169754 124856 169760 124908
rect 169812 124896 169818 124908
rect 261018 124896 261024 124908
rect 169812 124868 261024 124896
rect 169812 124856 169818 124868
rect 261018 124856 261024 124868
rect 261076 124856 261082 124908
rect 269850 124856 269856 124908
rect 269908 124896 269914 124908
rect 277578 124896 277584 124908
rect 269908 124868 277584 124896
rect 269908 124856 269914 124868
rect 277578 124856 277584 124868
rect 277636 124856 277642 124908
rect 296070 124856 296076 124908
rect 296128 124896 296134 124908
rect 354674 124896 354680 124908
rect 296128 124868 354680 124896
rect 296128 124856 296134 124868
rect 354674 124856 354680 124868
rect 354732 124856 354738 124908
rect 278130 124448 278136 124500
rect 278188 124488 278194 124500
rect 280246 124488 280252 124500
rect 278188 124460 280252 124488
rect 278188 124448 278194 124460
rect 280246 124448 280252 124460
rect 280304 124448 280310 124500
rect 226334 123496 226340 123548
rect 226392 123536 226398 123548
rect 270678 123536 270684 123548
rect 226392 123508 270684 123536
rect 226392 123496 226398 123508
rect 270678 123496 270684 123508
rect 270736 123496 270742 123548
rect 158714 123428 158720 123480
rect 158772 123468 158778 123480
rect 258166 123468 258172 123480
rect 158772 123440 258172 123468
rect 158772 123428 158778 123440
rect 258166 123428 258172 123440
rect 258224 123428 258230 123480
rect 133874 122068 133880 122120
rect 133932 122108 133938 122120
rect 254026 122108 254032 122120
rect 133932 122080 254032 122108
rect 133932 122068 133938 122080
rect 254026 122068 254032 122080
rect 254084 122068 254090 122120
rect 254578 122068 254584 122120
rect 254636 122108 254642 122120
rect 274818 122108 274824 122120
rect 254636 122080 274824 122108
rect 254636 122068 254642 122080
rect 274818 122068 274824 122080
rect 274876 122068 274882 122120
rect 136634 120708 136640 120760
rect 136692 120748 136698 120760
rect 255590 120748 255596 120760
rect 136692 120720 255596 120748
rect 136692 120708 136698 120720
rect 255590 120708 255596 120720
rect 255648 120708 255654 120760
rect 140774 119348 140780 119400
rect 140832 119388 140838 119400
rect 255498 119388 255504 119400
rect 140832 119360 255504 119388
rect 140832 119348 140838 119360
rect 255498 119348 255504 119360
rect 255556 119348 255562 119400
rect 151906 117920 151912 117972
rect 151964 117960 151970 117972
rect 256786 117960 256792 117972
rect 151964 117932 256792 117960
rect 151964 117920 151970 117932
rect 256786 117920 256792 117932
rect 256844 117920 256850 117972
rect 143626 116560 143632 116612
rect 143684 116600 143690 116612
rect 255406 116600 255412 116612
rect 143684 116572 255412 116600
rect 143684 116560 143690 116572
rect 255406 116560 255412 116572
rect 255464 116560 255470 116612
rect 127066 115200 127072 115252
rect 127124 115240 127130 115252
rect 252922 115240 252928 115252
rect 127124 115212 252928 115240
rect 127124 115200 127130 115212
rect 252922 115200 252928 115212
rect 252980 115200 252986 115252
rect 162854 113772 162860 113824
rect 162912 113812 162918 113824
rect 259638 113812 259644 113824
rect 162912 113784 259644 113812
rect 162912 113772 162918 113784
rect 259638 113772 259644 113784
rect 259696 113772 259702 113824
rect 460198 113092 460204 113144
rect 460256 113132 460262 113144
rect 579798 113132 579804 113144
rect 460256 113104 579804 113132
rect 460256 113092 460262 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 166994 112412 167000 112464
rect 167052 112452 167058 112464
rect 259546 112452 259552 112464
rect 167052 112424 259552 112452
rect 167052 112412 167058 112424
rect 259546 112412 259552 112424
rect 259604 112412 259610 112464
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 82078 111772 82084 111784
rect 3200 111744 82084 111772
rect 3200 111732 3206 111744
rect 82078 111732 82084 111744
rect 82136 111732 82142 111784
rect 173894 111052 173900 111104
rect 173952 111092 173958 111104
rect 260926 111092 260932 111104
rect 173952 111064 260932 111092
rect 173952 111052 173958 111064
rect 260926 111052 260932 111064
rect 260984 111052 260990 111104
rect 180794 109692 180800 109744
rect 180852 109732 180858 109744
rect 262306 109732 262312 109744
rect 180852 109704 262312 109732
rect 180852 109692 180858 109704
rect 262306 109692 262312 109704
rect 262364 109692 262370 109744
rect 185026 108264 185032 108316
rect 185084 108304 185090 108316
rect 263686 108304 263692 108316
rect 185084 108276 263692 108304
rect 185084 108264 185090 108276
rect 263686 108264 263692 108276
rect 263744 108264 263750 108316
rect 198734 106904 198740 106956
rect 198792 106944 198798 106956
rect 266446 106944 266452 106956
rect 198792 106916 266452 106944
rect 198792 106904 198798 106916
rect 266446 106904 266452 106916
rect 266504 106904 266510 106956
rect 187694 105544 187700 105596
rect 187752 105584 187758 105596
rect 263594 105584 263600 105596
rect 187752 105556 263600 105584
rect 187752 105544 187758 105556
rect 263594 105544 263600 105556
rect 263652 105544 263658 105596
rect 205634 104116 205640 104168
rect 205692 104156 205698 104168
rect 267826 104156 267832 104168
rect 205692 104128 267832 104156
rect 205692 104116 205698 104128
rect 267826 104116 267832 104128
rect 267884 104116 267890 104168
rect 223574 102824 223580 102876
rect 223632 102864 223638 102876
rect 270586 102864 270592 102876
rect 223632 102836 270592 102864
rect 223632 102824 223638 102836
rect 270586 102824 270592 102836
rect 270644 102824 270650 102876
rect 118694 102756 118700 102808
rect 118752 102796 118758 102808
rect 251450 102796 251456 102808
rect 118752 102768 251456 102796
rect 118752 102756 118758 102768
rect 251450 102756 251456 102768
rect 251508 102756 251514 102808
rect 135346 101396 135352 101448
rect 135404 101436 135410 101448
rect 254394 101436 254400 101448
rect 135404 101408 254400 101436
rect 135404 101396 135410 101408
rect 254394 101396 254400 101408
rect 254452 101396 254458 101448
rect 234706 99968 234712 100020
rect 234764 100008 234770 100020
rect 272334 100008 272340 100020
rect 234764 99980 272340 100008
rect 234764 99968 234770 99980
rect 272334 99968 272340 99980
rect 272392 99968 272398 100020
rect 144914 98608 144920 98660
rect 144972 98648 144978 98660
rect 256694 98648 256700 98660
rect 144972 98620 256700 98648
rect 144972 98608 144978 98620
rect 256694 98608 256700 98620
rect 256752 98608 256758 98660
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 57238 97968 57244 97980
rect 3568 97940 57244 97968
rect 3568 97928 3574 97940
rect 57238 97928 57244 97940
rect 57296 97928 57302 97980
rect 155954 97248 155960 97300
rect 156012 97288 156018 97300
rect 258534 97288 258540 97300
rect 156012 97260 258540 97288
rect 156012 97248 156018 97260
rect 258534 97248 258540 97260
rect 258592 97248 258598 97300
rect 111794 94460 111800 94512
rect 111852 94500 111858 94512
rect 249886 94500 249892 94512
rect 111852 94472 249892 94500
rect 111852 94460 111858 94472
rect 249886 94460 249892 94472
rect 249944 94460 249950 94512
rect 115934 93100 115940 93152
rect 115992 93140 115998 93152
rect 251358 93140 251364 93152
rect 115992 93112 251364 93140
rect 115992 93100 115998 93112
rect 251358 93100 251364 93112
rect 251416 93100 251422 93152
rect 106274 91740 106280 91792
rect 106332 91780 106338 91792
rect 248598 91780 248604 91792
rect 106332 91752 248604 91780
rect 106332 91740 106338 91752
rect 248598 91740 248604 91752
rect 248656 91740 248662 91792
rect 99374 90312 99380 90364
rect 99432 90352 99438 90364
rect 247402 90352 247408 90364
rect 99432 90324 247408 90352
rect 99432 90312 99438 90324
rect 247402 90312 247408 90324
rect 247460 90312 247466 90364
rect 49694 88952 49700 89004
rect 49752 88992 49758 89004
rect 239214 88992 239220 89004
rect 49752 88964 239220 88992
rect 49752 88952 49758 88964
rect 239214 88952 239220 88964
rect 239272 88952 239278 89004
rect 117314 87592 117320 87644
rect 117372 87632 117378 87644
rect 251266 87632 251272 87644
rect 117372 87604 251272 87632
rect 117372 87592 117378 87604
rect 251266 87592 251272 87604
rect 251324 87592 251330 87644
rect 113174 86232 113180 86284
rect 113232 86272 113238 86284
rect 250070 86272 250076 86284
rect 113232 86244 250076 86272
rect 113232 86232 113238 86244
rect 250070 86232 250076 86244
rect 250128 86232 250134 86284
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 79318 85524 79324 85536
rect 3568 85496 79324 85524
rect 3568 85484 3574 85496
rect 79318 85484 79324 85496
rect 79376 85484 79382 85536
rect 446398 73108 446404 73160
rect 446456 73148 446462 73160
rect 580166 73148 580172 73160
rect 446456 73120 580172 73148
rect 446456 73108 446462 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 142154 54476 142160 54528
rect 142212 54516 142218 54528
rect 255866 54516 255872 54528
rect 142212 54488 255872 54516
rect 142212 54476 142218 54488
rect 255866 54476 255872 54488
rect 255924 54476 255930 54528
rect 194594 53048 194600 53100
rect 194652 53088 194658 53100
rect 264974 53088 264980 53100
rect 194652 53060 264980 53088
rect 194652 53048 194658 53060
rect 264974 53048 264980 53060
rect 265032 53048 265038 53100
rect 494698 33056 494704 33108
rect 494756 33096 494762 33108
rect 580166 33096 580172 33108
rect 494756 33068 580172 33096
rect 494756 33056 494762 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 47578 32376 47584 32428
rect 47636 32416 47642 32428
rect 237742 32416 237748 32428
rect 47636 32388 237748 32416
rect 47636 32376 47642 32388
rect 237742 32376 237748 32388
rect 237800 32376 237806 32428
rect 295978 29588 295984 29640
rect 296036 29628 296042 29640
rect 347774 29628 347780 29640
rect 296036 29600 347780 29628
rect 296036 29588 296042 29600
rect 347774 29588 347780 29600
rect 347832 29588 347838 29640
rect 110506 24080 110512 24132
rect 110564 24120 110570 24132
rect 246390 24120 246396 24132
rect 110564 24092 246396 24120
rect 110564 24080 110570 24092
rect 246390 24080 246396 24092
rect 246448 24080 246454 24132
rect 102134 22720 102140 22772
rect 102192 22760 102198 22772
rect 246298 22760 246304 22772
rect 102192 22732 246304 22760
rect 102192 22720 102198 22732
rect 246298 22720 246304 22732
rect 246356 22720 246362 22772
rect 212534 21360 212540 21412
rect 212592 21400 212598 21412
rect 269114 21400 269120 21412
rect 212592 21372 269120 21400
rect 212592 21360 212598 21372
rect 269114 21360 269120 21372
rect 269172 21360 269178 21412
rect 209866 19932 209872 19984
rect 209924 19972 209930 19984
rect 267734 19972 267740 19984
rect 209924 19944 267740 19972
rect 209924 19932 209930 19944
rect 267734 19932 267740 19944
rect 267792 19932 267798 19984
rect 201586 18572 201592 18624
rect 201644 18612 201650 18624
rect 266906 18612 266912 18624
rect 201644 18584 266912 18612
rect 201644 18572 201650 18584
rect 266906 18572 266912 18584
rect 266964 18572 266970 18624
rect 160186 17280 160192 17332
rect 160244 17320 160250 17332
rect 260006 17320 260012 17332
rect 160244 17292 260012 17320
rect 160244 17280 160250 17292
rect 260006 17280 260012 17292
rect 260064 17280 260070 17332
rect 259546 17212 259552 17264
rect 259604 17252 259610 17264
rect 277486 17252 277492 17264
rect 259604 17224 277492 17252
rect 259604 17212 259610 17224
rect 277486 17212 277492 17224
rect 277544 17212 277550 17264
rect 292574 17212 292580 17264
rect 292632 17252 292638 17264
rect 343634 17252 343640 17264
rect 292632 17224 343640 17252
rect 292632 17212 292638 17224
rect 343634 17212 343640 17224
rect 343692 17212 343698 17264
rect 177850 15852 177856 15904
rect 177908 15892 177914 15904
rect 262674 15892 262680 15904
rect 177908 15864 262680 15892
rect 177908 15852 177914 15864
rect 262674 15852 262680 15864
rect 262732 15852 262738 15904
rect 289814 15852 289820 15904
rect 289872 15892 289878 15904
rect 330386 15892 330392 15904
rect 289872 15864 330392 15892
rect 289872 15852 289878 15864
rect 330386 15852 330392 15864
rect 330444 15852 330450 15904
rect 120626 14424 120632 14476
rect 120684 14464 120690 14476
rect 247678 14464 247684 14476
rect 120684 14436 247684 14464
rect 120684 14424 120690 14436
rect 247678 14424 247684 14436
rect 247736 14424 247742 14476
rect 264146 14424 264152 14476
rect 264204 14464 264210 14476
rect 277394 14464 277400 14476
rect 264204 14436 277400 14464
rect 264204 14424 264210 14436
rect 277394 14424 277400 14436
rect 277452 14424 277458 14476
rect 287146 14424 287152 14476
rect 287204 14464 287210 14476
rect 312170 14464 312176 14476
rect 287204 14436 312176 14464
rect 287204 14424 287210 14436
rect 312170 14424 312176 14436
rect 312228 14424 312234 14476
rect 260190 13132 260196 13184
rect 260248 13172 260254 13184
rect 276106 13172 276112 13184
rect 260248 13144 276112 13172
rect 260248 13132 260254 13144
rect 276106 13132 276112 13144
rect 276164 13132 276170 13184
rect 123018 13064 123024 13116
rect 123076 13104 123082 13116
rect 250438 13104 250444 13116
rect 123076 13076 250444 13104
rect 123076 13064 123082 13076
rect 250438 13064 250444 13076
rect 250496 13064 250502 13116
rect 276014 13064 276020 13116
rect 276072 13104 276078 13116
rect 280522 13104 280528 13116
rect 276072 13076 280528 13104
rect 276072 13064 276078 13076
rect 280522 13064 280528 13076
rect 280580 13064 280586 13116
rect 285674 13064 285680 13116
rect 285732 13104 285738 13116
rect 307938 13104 307944 13116
rect 285732 13076 307944 13104
rect 285732 13064 285738 13076
rect 307938 13064 307944 13076
rect 307996 13064 308002 13116
rect 255866 12452 255872 12504
rect 255924 12492 255930 12504
rect 257338 12492 257344 12504
rect 255924 12464 257344 12492
rect 255924 12452 255930 12464
rect 257338 12452 257344 12464
rect 257396 12452 257402 12504
rect 160094 11772 160100 11824
rect 160152 11812 160158 11824
rect 161290 11812 161296 11824
rect 160152 11784 161296 11812
rect 160152 11772 160158 11784
rect 161290 11772 161296 11784
rect 161348 11772 161354 11824
rect 184934 11772 184940 11824
rect 184992 11812 184998 11824
rect 186130 11812 186136 11824
rect 184992 11784 186136 11812
rect 184992 11772 184998 11784
rect 186130 11772 186136 11784
rect 186188 11772 186194 11824
rect 234614 11772 234620 11824
rect 234672 11812 234678 11824
rect 235810 11812 235816 11824
rect 234672 11784 235816 11812
rect 234672 11772 234678 11784
rect 235810 11772 235816 11784
rect 235868 11772 235874 11824
rect 284938 11772 284944 11824
rect 284996 11812 285002 11824
rect 293218 11812 293224 11824
rect 284996 11784 293224 11812
rect 284996 11772 285002 11784
rect 293218 11772 293224 11784
rect 293276 11772 293282 11824
rect 105722 11704 105728 11756
rect 105780 11744 105786 11756
rect 248506 11744 248512 11756
rect 105780 11716 248512 11744
rect 105780 11704 105786 11716
rect 248506 11704 248512 11716
rect 248564 11704 248570 11756
rect 266538 11704 266544 11756
rect 266596 11744 266602 11756
rect 278038 11744 278044 11756
rect 266596 11716 278044 11744
rect 266596 11704 266602 11716
rect 278038 11704 278044 11716
rect 278096 11704 278102 11756
rect 287054 11704 287060 11756
rect 287112 11744 287118 11756
rect 316218 11744 316224 11756
rect 287112 11716 316224 11744
rect 287112 11704 287118 11716
rect 316218 11704 316224 11716
rect 316276 11704 316282 11756
rect 272426 10480 272432 10532
rect 272484 10520 272490 10532
rect 279326 10520 279332 10532
rect 272484 10492 279332 10520
rect 272484 10480 272490 10492
rect 279326 10480 279332 10492
rect 279384 10480 279390 10532
rect 60826 10276 60832 10328
rect 60884 10316 60890 10328
rect 239398 10316 239404 10328
rect 60884 10288 239404 10316
rect 60884 10276 60890 10288
rect 239398 10276 239404 10288
rect 239456 10276 239462 10328
rect 244642 10276 244648 10328
rect 244700 10316 244706 10328
rect 274726 10316 274732 10328
rect 244700 10288 274732 10316
rect 244700 10276 244706 10288
rect 274726 10276 274732 10288
rect 274784 10276 274790 10328
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 241698 8984 241704 9036
rect 241756 9024 241762 9036
rect 273438 9024 273444 9036
rect 241756 8996 273444 9024
rect 241756 8984 241762 8996
rect 273438 8984 273444 8996
rect 273496 8984 273502 9036
rect 109310 8916 109316 8968
rect 109368 8956 109374 8968
rect 243538 8956 243544 8968
rect 109368 8928 243544 8956
rect 109368 8916 109374 8928
rect 243538 8916 243544 8928
rect 243596 8916 243602 8968
rect 299014 8916 299020 8968
rect 299072 8956 299078 8968
rect 401318 8956 401324 8968
rect 299072 8928 401324 8956
rect 299072 8916 299078 8928
rect 401318 8916 401324 8928
rect 401376 8916 401382 8968
rect 271230 8236 271236 8288
rect 271288 8276 271294 8288
rect 275278 8276 275284 8288
rect 271288 8248 275284 8276
rect 271288 8236 271294 8248
rect 275278 8236 275284 8248
rect 275336 8236 275342 8288
rect 248782 7624 248788 7676
rect 248840 7664 248846 7676
rect 268378 7664 268384 7676
rect 248840 7636 268384 7664
rect 248840 7624 248846 7636
rect 268378 7624 268384 7636
rect 268436 7624 268442 7676
rect 70302 7556 70308 7608
rect 70360 7596 70366 7608
rect 242158 7596 242164 7608
rect 70360 7568 242164 7596
rect 70360 7556 70366 7568
rect 242158 7556 242164 7568
rect 242216 7556 242222 7608
rect 247586 7556 247592 7608
rect 247644 7596 247650 7608
rect 275094 7596 275100 7608
rect 247644 7568 275100 7596
rect 247644 7556 247650 7568
rect 275094 7556 275100 7568
rect 275152 7556 275158 7608
rect 298094 7556 298100 7608
rect 298152 7596 298158 7608
rect 372890 7596 372896 7608
rect 298152 7568 372896 7596
rect 298152 7556 298158 7568
rect 372890 7556 372896 7568
rect 372948 7556 372954 7608
rect 283098 6876 283104 6928
rect 283156 6916 283162 6928
rect 288986 6916 288992 6928
rect 283156 6888 288992 6916
rect 283156 6876 283162 6888
rect 288986 6876 288992 6888
rect 289044 6876 289050 6928
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 44818 6848 44824 6860
rect 3476 6820 44824 6848
rect 3476 6808 3482 6820
rect 44818 6808 44824 6820
rect 44876 6808 44882 6860
rect 289078 6808 289084 6860
rect 289136 6848 289142 6860
rect 309042 6848 309048 6860
rect 289136 6820 309048 6848
rect 289136 6808 289142 6820
rect 309042 6808 309048 6820
rect 309100 6808 309106 6860
rect 283006 6740 283012 6792
rect 283064 6780 283070 6792
rect 294874 6780 294880 6792
rect 283064 6752 294880 6780
rect 283064 6740 283070 6752
rect 294874 6740 294880 6752
rect 294932 6740 294938 6792
rect 295518 6740 295524 6792
rect 295576 6780 295582 6792
rect 358722 6780 358728 6792
rect 295576 6752 358728 6780
rect 295576 6740 295582 6752
rect 358722 6740 358728 6752
rect 358780 6740 358786 6792
rect 292482 6672 292488 6724
rect 292540 6712 292546 6724
rect 382366 6712 382372 6724
rect 292540 6684 382372 6712
rect 292540 6672 292546 6684
rect 382366 6672 382372 6684
rect 382424 6672 382430 6724
rect 291010 6604 291016 6656
rect 291068 6644 291074 6656
rect 385954 6644 385960 6656
rect 291068 6616 385960 6644
rect 291068 6604 291074 6616
rect 385954 6604 385960 6616
rect 386012 6604 386018 6656
rect 289262 6536 289268 6588
rect 289320 6576 289326 6588
rect 396534 6576 396540 6588
rect 289320 6548 396540 6576
rect 289320 6536 289326 6548
rect 396534 6536 396540 6548
rect 396592 6536 396598 6588
rect 289630 6468 289636 6520
rect 289688 6508 289694 6520
rect 400122 6508 400128 6520
rect 289688 6480 400128 6508
rect 289688 6468 289694 6480
rect 400122 6468 400128 6480
rect 400180 6468 400186 6520
rect 289446 6400 289452 6452
rect 289504 6440 289510 6452
rect 403618 6440 403624 6452
rect 289504 6412 403624 6440
rect 289504 6400 289510 6412
rect 403618 6400 403624 6412
rect 403676 6400 403682 6452
rect 289354 6332 289360 6384
rect 289412 6372 289418 6384
rect 407206 6372 407212 6384
rect 289412 6344 407212 6372
rect 289412 6332 289418 6344
rect 407206 6332 407212 6344
rect 407264 6332 407270 6384
rect 290918 6264 290924 6316
rect 290976 6304 290982 6316
rect 410794 6304 410800 6316
rect 290976 6276 410800 6304
rect 290976 6264 290982 6276
rect 410794 6264 410800 6276
rect 410852 6264 410858 6316
rect 238110 6196 238116 6248
rect 238168 6236 238174 6248
rect 273346 6236 273352 6248
rect 238168 6208 273352 6236
rect 238168 6196 238174 6208
rect 273346 6196 273352 6208
rect 273404 6196 273410 6248
rect 290734 6196 290740 6248
rect 290792 6236 290798 6248
rect 416682 6236 416688 6248
rect 290792 6208 416688 6236
rect 290792 6196 290798 6208
rect 416682 6196 416688 6208
rect 416740 6196 416746 6248
rect 119890 6128 119896 6180
rect 119948 6168 119954 6180
rect 251634 6168 251640 6180
rect 119948 6140 251640 6168
rect 119948 6128 119954 6140
rect 251634 6128 251640 6140
rect 251692 6128 251698 6180
rect 254670 6128 254676 6180
rect 254728 6168 254734 6180
rect 276474 6168 276480 6180
rect 254728 6140 276480 6168
rect 254728 6128 254734 6140
rect 276474 6128 276480 6140
rect 276532 6128 276538 6180
rect 292390 6128 292396 6180
rect 292448 6168 292454 6180
rect 420178 6168 420184 6180
rect 292448 6140 420184 6168
rect 292448 6128 292454 6140
rect 420178 6128 420184 6140
rect 420236 6128 420242 6180
rect 281810 5516 281816 5568
rect 281868 5556 281874 5568
rect 284202 5556 284208 5568
rect 281868 5528 284208 5556
rect 281868 5516 281874 5528
rect 284202 5516 284208 5528
rect 284260 5516 284266 5568
rect 240502 4904 240508 4956
rect 240560 4944 240566 4956
rect 273254 4944 273260 4956
rect 240560 4916 273260 4944
rect 240560 4904 240566 4916
rect 273254 4904 273260 4916
rect 273312 4904 273318 4956
rect 283466 4904 283472 4956
rect 283524 4944 283530 4956
rect 290182 4944 290188 4956
rect 283524 4916 290188 4944
rect 283524 4904 283530 4916
rect 290182 4904 290188 4916
rect 290240 4904 290246 4956
rect 227530 4836 227536 4888
rect 227588 4876 227594 4888
rect 270494 4876 270500 4888
rect 227588 4848 270500 4876
rect 227588 4836 227594 4848
rect 270494 4836 270500 4848
rect 270552 4836 270558 4888
rect 286318 4836 286324 4888
rect 286376 4876 286382 4888
rect 297266 4876 297272 4888
rect 286376 4848 297272 4876
rect 286376 4836 286382 4848
rect 297266 4836 297272 4848
rect 297324 4836 297330 4888
rect 80882 4768 80888 4820
rect 80940 4808 80946 4820
rect 244550 4808 244556 4820
rect 80940 4780 244556 4808
rect 80940 4768 80946 4780
rect 244550 4768 244556 4780
rect 244608 4768 244614 4820
rect 284294 4768 284300 4820
rect 284352 4808 284358 4820
rect 298462 4808 298468 4820
rect 284352 4780 298468 4808
rect 284352 4768 284358 4780
rect 298462 4768 298468 4780
rect 298520 4768 298526 4820
rect 278314 4156 278320 4208
rect 278372 4196 278378 4208
rect 279418 4196 279424 4208
rect 278372 4168 279424 4196
rect 278372 4156 278378 4168
rect 279418 4156 279424 4168
rect 279476 4156 279482 4208
rect 281718 4156 281724 4208
rect 281776 4196 281782 4208
rect 285398 4196 285404 4208
rect 281776 4168 285404 4196
rect 281776 4156 281782 4168
rect 285398 4156 285404 4168
rect 285456 4156 285462 4208
rect 299566 4156 299572 4208
rect 299624 4196 299630 4208
rect 300762 4196 300768 4208
rect 299624 4168 300768 4196
rect 299624 4156 299630 4168
rect 300762 4156 300768 4168
rect 300820 4156 300826 4208
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 7558 4128 7564 4140
rect 2924 4100 7564 4128
rect 2924 4088 2930 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 45462 4088 45468 4140
rect 45520 4128 45526 4140
rect 46290 4128 46296 4140
rect 45520 4100 46296 4128
rect 45520 4088 45526 4100
rect 46290 4088 46296 4100
rect 46348 4088 46354 4140
rect 257062 4088 257068 4140
rect 257120 4128 257126 4140
rect 260190 4128 260196 4140
rect 257120 4100 260196 4128
rect 257120 4088 257126 4100
rect 260190 4088 260196 4100
rect 260248 4088 260254 4140
rect 277118 4088 277124 4140
rect 277176 4128 277182 4140
rect 279510 4128 279516 4140
rect 277176 4100 279516 4128
rect 277176 4088 277182 4100
rect 279510 4088 279516 4100
rect 279568 4088 279574 4140
rect 288342 4088 288348 4140
rect 288400 4128 288406 4140
rect 335078 4128 335084 4140
rect 288400 4100 335084 4128
rect 288400 4088 288406 4100
rect 335078 4088 335084 4100
rect 335136 4088 335142 4140
rect 338758 4088 338764 4140
rect 338816 4128 338822 4140
rect 371694 4128 371700 4140
rect 338816 4100 371700 4128
rect 338816 4088 338822 4100
rect 371694 4088 371700 4100
rect 371752 4088 371758 4140
rect 434438 4088 434444 4140
rect 434496 4128 434502 4140
rect 439130 4128 439136 4140
rect 434496 4100 439136 4128
rect 434496 4088 434502 4100
rect 439130 4088 439136 4100
rect 439188 4088 439194 4140
rect 536190 4088 536196 4140
rect 536248 4128 536254 4140
rect 538398 4128 538404 4140
rect 536248 4100 538404 4128
rect 536248 4088 536254 4100
rect 538398 4088 538404 4100
rect 538456 4088 538462 4140
rect 295334 4020 295340 4072
rect 295392 4060 295398 4072
rect 356330 4060 356336 4072
rect 295392 4032 356336 4060
rect 295392 4020 295398 4032
rect 356330 4020 356336 4032
rect 356388 4020 356394 4072
rect 428458 4020 428464 4072
rect 428516 4060 428522 4072
rect 439406 4060 439412 4072
rect 428516 4032 439412 4060
rect 428516 4020 428522 4032
rect 439406 4020 439412 4032
rect 439464 4020 439470 4072
rect 246390 3952 246396 4004
rect 246448 3992 246454 4004
rect 253290 3992 253296 4004
rect 246448 3964 253296 3992
rect 246448 3952 246454 3964
rect 253290 3952 253296 3964
rect 253348 3952 253354 4004
rect 295426 3952 295432 4004
rect 295484 3992 295490 4004
rect 359918 3992 359924 4004
rect 295484 3964 359924 3992
rect 295484 3952 295490 3964
rect 359918 3952 359924 3964
rect 359976 3952 359982 4004
rect 427262 3952 427268 4004
rect 427320 3992 427326 4004
rect 439222 3992 439228 4004
rect 427320 3964 439228 3992
rect 427320 3952 427326 3964
rect 439222 3952 439228 3964
rect 439280 3952 439286 4004
rect 244090 3884 244096 3936
rect 244148 3924 244154 3936
rect 254578 3924 254584 3936
rect 244148 3896 254584 3924
rect 244148 3884 244154 3896
rect 254578 3884 254584 3896
rect 254636 3884 254642 3936
rect 295242 3884 295248 3936
rect 295300 3924 295306 3936
rect 381170 3924 381176 3936
rect 295300 3896 381176 3924
rect 295300 3884 295306 3896
rect 381170 3884 381176 3896
rect 381228 3884 381234 3936
rect 426158 3884 426164 3936
rect 426216 3924 426222 3936
rect 438854 3924 438860 3936
rect 426216 3896 438860 3924
rect 426216 3884 426222 3896
rect 438854 3884 438860 3896
rect 438912 3884 438918 3936
rect 239306 3816 239312 3868
rect 239364 3856 239370 3868
rect 253382 3856 253388 3868
rect 239364 3828 253388 3856
rect 239364 3816 239370 3828
rect 253382 3816 253388 3828
rect 253440 3816 253446 3868
rect 258166 3816 258172 3868
rect 258224 3856 258230 3868
rect 265618 3856 265624 3868
rect 258224 3828 265624 3856
rect 258224 3816 258230 3828
rect 265618 3816 265624 3828
rect 265676 3816 265682 3868
rect 291102 3816 291108 3868
rect 291160 3856 291166 3868
rect 378870 3856 378876 3868
rect 291160 3828 378876 3856
rect 291160 3816 291166 3828
rect 378870 3816 378876 3828
rect 378928 3816 378934 3868
rect 424962 3816 424968 3868
rect 425020 3856 425026 3868
rect 437658 3856 437664 3868
rect 425020 3828 437664 3856
rect 425020 3816 425026 3828
rect 437658 3816 437664 3828
rect 437716 3816 437722 3868
rect 516778 3816 516784 3868
rect 516836 3856 516842 3868
rect 519538 3856 519544 3868
rect 516836 3828 519544 3856
rect 516836 3816 516842 3828
rect 519538 3816 519544 3828
rect 519596 3816 519602 3868
rect 574738 3816 574744 3868
rect 574796 3856 574802 3868
rect 577406 3856 577412 3868
rect 574796 3828 577412 3856
rect 574796 3816 574802 3828
rect 577406 3816 577412 3828
rect 577464 3816 577470 3868
rect 35986 3748 35992 3800
rect 36044 3788 36050 3800
rect 46198 3788 46204 3800
rect 36044 3760 46204 3788
rect 36044 3748 36050 3760
rect 46198 3748 46204 3760
rect 46256 3748 46262 3800
rect 135254 3748 135260 3800
rect 135312 3788 135318 3800
rect 136450 3788 136456 3800
rect 135312 3760 136456 3788
rect 135312 3748 135318 3760
rect 136450 3748 136456 3760
rect 136508 3748 136514 3800
rect 171962 3748 171968 3800
rect 172020 3788 172026 3800
rect 261386 3788 261392 3800
rect 172020 3760 261392 3788
rect 172020 3748 172026 3760
rect 261386 3748 261392 3760
rect 261444 3748 261450 3800
rect 295150 3748 295156 3800
rect 295208 3788 295214 3800
rect 388254 3788 388260 3800
rect 295208 3760 388260 3788
rect 295208 3748 295214 3760
rect 388254 3748 388260 3760
rect 388312 3748 388318 3800
rect 423766 3748 423772 3800
rect 423824 3788 423830 3800
rect 437842 3788 437848 3800
rect 423824 3760 437848 3788
rect 423824 3748 423830 3760
rect 437842 3748 437848 3760
rect 437900 3748 437906 3800
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 39298 3720 39304 3732
rect 11204 3692 39304 3720
rect 11204 3680 11210 3692
rect 39298 3680 39304 3692
rect 39356 3680 39362 3732
rect 53742 3680 53748 3732
rect 53800 3720 53806 3732
rect 54478 3720 54484 3732
rect 53800 3692 54484 3720
rect 53800 3680 53806 3692
rect 54478 3680 54484 3692
rect 54536 3680 54542 3732
rect 82078 3680 82084 3732
rect 82136 3720 82142 3732
rect 93118 3720 93124 3732
rect 82136 3692 93124 3720
rect 82136 3680 82142 3692
rect 93118 3680 93124 3692
rect 93176 3680 93182 3732
rect 124674 3680 124680 3732
rect 124732 3720 124738 3732
rect 238018 3720 238024 3732
rect 124732 3692 238024 3720
rect 124732 3680 124738 3692
rect 238018 3680 238024 3692
rect 238076 3680 238082 3732
rect 242894 3680 242900 3732
rect 242952 3720 242958 3732
rect 264238 3720 264244 3732
rect 242952 3692 264244 3720
rect 242952 3680 242958 3692
rect 264238 3680 264244 3692
rect 264296 3680 264302 3732
rect 289722 3680 289728 3732
rect 289780 3720 289786 3732
rect 395338 3720 395344 3732
rect 289780 3692 395344 3720
rect 289780 3680 289786 3692
rect 395338 3680 395344 3692
rect 395396 3680 395402 3732
rect 422570 3680 422576 3732
rect 422628 3720 422634 3732
rect 437474 3720 437480 3732
rect 422628 3692 437480 3720
rect 422628 3680 422634 3692
rect 437474 3680 437480 3692
rect 437532 3680 437538 3732
rect 462958 3680 462964 3732
rect 463016 3720 463022 3732
rect 463016 3692 470594 3720
rect 463016 3680 463022 3692
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 95878 3652 95884 3664
rect 39632 3624 95884 3652
rect 39632 3612 39638 3624
rect 95878 3612 95884 3624
rect 95936 3612 95942 3664
rect 96246 3612 96252 3664
rect 96304 3652 96310 3664
rect 97258 3652 97264 3664
rect 96304 3624 97264 3652
rect 96304 3612 96310 3624
rect 97258 3612 97264 3624
rect 97316 3612 97322 3664
rect 102226 3612 102232 3664
rect 102284 3652 102290 3664
rect 248690 3652 248696 3664
rect 102284 3624 248696 3652
rect 102284 3612 102290 3624
rect 248690 3612 248696 3624
rect 248748 3612 248754 3664
rect 251174 3612 251180 3664
rect 251232 3652 251238 3664
rect 261478 3652 261484 3664
rect 251232 3624 261484 3652
rect 251232 3612 251238 3624
rect 261478 3612 261484 3624
rect 261536 3612 261542 3664
rect 293494 3612 293500 3664
rect 293552 3652 293558 3664
rect 402514 3652 402520 3664
rect 293552 3624 402520 3652
rect 293552 3612 293558 3624
rect 402514 3612 402520 3624
rect 402572 3612 402578 3664
rect 421374 3612 421380 3664
rect 421432 3652 421438 3664
rect 439038 3652 439044 3664
rect 421432 3624 439044 3652
rect 421432 3612 421438 3624
rect 439038 3612 439044 3624
rect 439096 3612 439102 3664
rect 442258 3612 442264 3664
rect 442316 3652 442322 3664
rect 447410 3652 447416 3664
rect 442316 3624 447416 3652
rect 442316 3612 442322 3624
rect 447410 3612 447416 3624
rect 447468 3612 447474 3664
rect 456058 3612 456064 3664
rect 456116 3652 456122 3664
rect 465166 3652 465172 3664
rect 456116 3624 465172 3652
rect 456116 3612 456122 3624
rect 465166 3612 465172 3624
rect 465224 3612 465230 3664
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 4798 3584 4804 3596
rect 1728 3556 4804 3584
rect 1728 3544 1734 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 10318 3584 10324 3596
rect 6886 3556 10324 3584
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 6886 3516 6914 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 13078 3584 13084 3596
rect 12400 3556 13084 3584
rect 12400 3544 12406 3556
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 21358 3584 21364 3596
rect 20680 3556 21364 3584
rect 20680 3544 20686 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 71038 3584 71044 3596
rect 25372 3556 71044 3584
rect 25372 3544 25378 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 71498 3544 71504 3596
rect 71556 3584 71562 3596
rect 72418 3584 72424 3596
rect 71556 3556 72424 3584
rect 71556 3544 71562 3556
rect 72418 3544 72424 3556
rect 72476 3544 72482 3596
rect 85666 3544 85672 3596
rect 85724 3584 85730 3596
rect 88978 3584 88984 3596
rect 85724 3556 88984 3584
rect 85724 3544 85730 3556
rect 88978 3544 88984 3556
rect 89036 3544 89042 3596
rect 89254 3544 89260 3596
rect 89312 3584 89318 3596
rect 244734 3584 244740 3596
rect 89312 3556 244740 3584
rect 89312 3544 89318 3556
rect 244734 3544 244740 3556
rect 244792 3544 244798 3596
rect 244826 3544 244832 3596
rect 244884 3544 244890 3596
rect 249978 3544 249984 3596
rect 250036 3584 250042 3596
rect 258166 3584 258172 3596
rect 250036 3556 258172 3584
rect 250036 3544 250042 3556
rect 258166 3544 258172 3556
rect 258224 3544 258230 3596
rect 258258 3544 258264 3596
rect 258316 3584 258322 3596
rect 260098 3584 260104 3596
rect 258316 3556 260104 3584
rect 258316 3544 258322 3556
rect 260098 3544 260104 3556
rect 260156 3544 260162 3596
rect 267734 3544 267740 3596
rect 267792 3584 267798 3596
rect 273898 3584 273904 3596
rect 267792 3556 273904 3584
rect 267792 3544 267798 3556
rect 273898 3544 273904 3556
rect 273956 3544 273962 3596
rect 281442 3544 281448 3596
rect 281500 3584 281506 3596
rect 281500 3556 287054 3584
rect 281500 3544 281506 3556
rect 4120 3488 6914 3516
rect 4120 3476 4126 3488
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8938 3516 8944 3528
rect 7708 3488 8944 3516
rect 7708 3476 7714 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 15988 3488 45554 3516
rect 15988 3476 15994 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 25498 3448 25504 3460
rect 624 3420 25504 3448
rect 624 3408 630 3420
rect 25498 3408 25504 3420
rect 25556 3408 25562 3460
rect 27706 3408 27712 3460
rect 27764 3448 27770 3460
rect 31018 3448 31024 3460
rect 27764 3420 31024 3448
rect 27764 3408 27770 3420
rect 31018 3408 31024 3420
rect 31076 3408 31082 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 35158 3448 35164 3460
rect 33652 3420 35164 3448
rect 33652 3408 33658 3420
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 38378 3408 38384 3460
rect 38436 3448 38442 3460
rect 39390 3448 39396 3460
rect 38436 3420 39396 3448
rect 38436 3408 38442 3420
rect 39390 3408 39396 3420
rect 39448 3408 39454 3460
rect 40678 3408 40684 3460
rect 40736 3448 40742 3460
rect 43438 3448 43444 3460
rect 40736 3420 43444 3448
rect 40736 3408 40742 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 45526 3448 45554 3488
rect 46658 3476 46664 3528
rect 46716 3516 46722 3528
rect 47578 3516 47584 3528
rect 46716 3488 47584 3516
rect 46716 3476 46722 3488
rect 47578 3476 47584 3488
rect 47636 3476 47642 3528
rect 47854 3476 47860 3528
rect 47912 3516 47918 3528
rect 48958 3516 48964 3528
rect 47912 3488 48964 3516
rect 47912 3476 47918 3488
rect 48958 3476 48964 3488
rect 49016 3476 49022 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 57330 3516 57336 3528
rect 56100 3488 57336 3516
rect 56100 3476 56106 3488
rect 57330 3476 57336 3488
rect 57388 3476 57394 3528
rect 60734 3476 60740 3528
rect 60792 3516 60798 3528
rect 61654 3516 61660 3528
rect 60792 3488 61660 3516
rect 60792 3476 60798 3488
rect 61654 3476 61660 3488
rect 61712 3476 61718 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 244844 3516 244872 3544
rect 83332 3488 244872 3516
rect 83332 3476 83338 3488
rect 253474 3476 253480 3528
rect 253532 3516 253538 3528
rect 269758 3516 269764 3528
rect 253532 3488 269764 3516
rect 253532 3476 253538 3488
rect 269758 3476 269764 3488
rect 269816 3476 269822 3528
rect 281626 3476 281632 3528
rect 281684 3516 281690 3528
rect 283098 3516 283104 3528
rect 281684 3488 283104 3516
rect 281684 3476 281690 3488
rect 283098 3476 283104 3488
rect 283156 3476 283162 3528
rect 287026 3516 287054 3556
rect 293862 3544 293868 3596
rect 293920 3584 293926 3596
rect 406010 3584 406016 3596
rect 293920 3556 406016 3584
rect 293920 3544 293926 3556
rect 406010 3544 406016 3556
rect 406068 3544 406074 3596
rect 418982 3544 418988 3596
rect 419040 3584 419046 3596
rect 438946 3584 438952 3596
rect 419040 3556 438952 3584
rect 419040 3544 419046 3556
rect 438946 3544 438952 3556
rect 439004 3544 439010 3596
rect 443638 3544 443644 3596
rect 443696 3584 443702 3596
rect 443696 3556 451274 3584
rect 443696 3544 443702 3556
rect 292574 3516 292580 3528
rect 287026 3488 292580 3516
rect 292574 3476 292580 3488
rect 292632 3476 292638 3528
rect 295058 3476 295064 3528
rect 295116 3516 295122 3528
rect 409598 3516 409604 3528
rect 295116 3488 409604 3516
rect 295116 3476 295122 3488
rect 409598 3476 409604 3488
rect 409656 3476 409662 3528
rect 417878 3476 417884 3528
rect 417936 3516 417942 3528
rect 437750 3516 437756 3528
rect 417936 3488 437756 3516
rect 417936 3476 417942 3488
rect 437750 3476 437756 3488
rect 437808 3476 437814 3528
rect 440234 3476 440240 3528
rect 440292 3516 440298 3528
rect 441522 3516 441528 3528
rect 440292 3488 441528 3516
rect 440292 3476 440298 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 448514 3476 448520 3528
rect 448572 3516 448578 3528
rect 449802 3516 449808 3528
rect 448572 3488 449808 3516
rect 448572 3476 448578 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 451246 3516 451274 3556
rect 453298 3544 453304 3596
rect 453356 3584 453362 3596
rect 455690 3584 455696 3596
rect 453356 3556 455696 3584
rect 453356 3544 453362 3556
rect 455690 3544 455696 3556
rect 455748 3544 455754 3596
rect 467098 3544 467104 3596
rect 467156 3584 467162 3596
rect 469858 3584 469864 3596
rect 467156 3556 469864 3584
rect 467156 3544 467162 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 470566 3584 470594 3692
rect 480530 3584 480536 3596
rect 470566 3556 480536 3584
rect 480530 3544 480536 3556
rect 480588 3544 480594 3596
rect 484026 3584 484032 3596
rect 481560 3556 484032 3584
rect 471054 3516 471060 3528
rect 451246 3488 471060 3516
rect 471054 3476 471060 3488
rect 471112 3476 471118 3528
rect 471238 3476 471244 3528
rect 471296 3516 471302 3528
rect 473446 3516 473452 3528
rect 471296 3488 473452 3516
rect 471296 3476 471302 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 476758 3476 476764 3528
rect 476816 3516 476822 3528
rect 481560 3516 481588 3556
rect 484026 3544 484032 3556
rect 484084 3544 484090 3596
rect 491938 3544 491944 3596
rect 491996 3584 492002 3596
rect 494698 3584 494704 3596
rect 491996 3556 494704 3584
rect 491996 3544 492002 3556
rect 494698 3544 494704 3556
rect 494756 3544 494762 3596
rect 500218 3544 500224 3596
rect 500276 3584 500282 3596
rect 501782 3584 501788 3596
rect 500276 3556 501788 3584
rect 500276 3544 500282 3556
rect 501782 3544 501788 3556
rect 501840 3544 501846 3596
rect 511258 3544 511264 3596
rect 511316 3584 511322 3596
rect 513558 3584 513564 3596
rect 511316 3556 513564 3584
rect 511316 3544 511322 3556
rect 513558 3544 513564 3556
rect 513616 3544 513622 3596
rect 514018 3544 514024 3596
rect 514076 3584 514082 3596
rect 515950 3584 515956 3596
rect 514076 3556 515956 3584
rect 514076 3544 514082 3556
rect 515950 3544 515956 3556
rect 516008 3544 516014 3596
rect 549898 3544 549904 3596
rect 549956 3584 549962 3596
rect 551462 3584 551468 3596
rect 549956 3556 551468 3584
rect 549956 3544 549962 3556
rect 551462 3544 551468 3556
rect 551520 3544 551526 3596
rect 476816 3488 481588 3516
rect 476816 3476 476822 3488
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 482462 3516 482468 3528
rect 481692 3488 482468 3516
rect 481692 3476 481698 3488
rect 482462 3476 482468 3488
rect 482520 3476 482526 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 496078 3476 496084 3528
rect 496136 3516 496142 3528
rect 497090 3516 497096 3528
rect 496136 3488 497096 3516
rect 496136 3476 496142 3488
rect 497090 3476 497096 3488
rect 497148 3476 497154 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 514110 3476 514116 3528
rect 514168 3516 514174 3528
rect 514754 3516 514760 3528
rect 514168 3488 514760 3516
rect 514168 3476 514174 3488
rect 514754 3476 514760 3488
rect 514812 3476 514818 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 523862 3516 523868 3528
rect 523092 3488 523868 3516
rect 523092 3476 523098 3488
rect 523862 3476 523868 3488
rect 523920 3476 523926 3528
rect 527910 3476 527916 3528
rect 527968 3516 527974 3528
rect 533706 3516 533712 3528
rect 527968 3488 533712 3516
rect 527968 3476 527974 3488
rect 533706 3476 533712 3488
rect 533764 3476 533770 3528
rect 547874 3476 547880 3528
rect 547932 3516 547938 3528
rect 548702 3516 548708 3528
rect 547932 3488 548708 3516
rect 547932 3476 547938 3488
rect 548702 3476 548708 3488
rect 548760 3476 548766 3528
rect 571978 3476 571984 3528
rect 572036 3516 572042 3528
rect 573910 3516 573916 3528
rect 572036 3488 573916 3516
rect 572036 3476 572042 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 580994 3476 581000 3528
rect 581052 3516 581058 3528
rect 581822 3516 581828 3528
rect 581052 3488 581828 3516
rect 581052 3476 581058 3488
rect 581822 3476 581828 3488
rect 581880 3476 581886 3528
rect 64138 3448 64144 3460
rect 45526 3420 64144 3448
rect 64138 3408 64144 3420
rect 64196 3408 64202 3460
rect 64322 3408 64328 3460
rect 64380 3448 64386 3460
rect 68278 3448 68284 3460
rect 64380 3420 68284 3448
rect 64380 3408 64386 3420
rect 68278 3408 68284 3420
rect 68336 3408 68342 3460
rect 79686 3408 79692 3460
rect 79744 3448 79750 3460
rect 244458 3448 244464 3460
rect 79744 3420 244464 3448
rect 79744 3408 79750 3420
rect 244458 3408 244464 3420
rect 244516 3408 244522 3460
rect 252370 3408 252376 3460
rect 252428 3448 252434 3460
rect 271138 3448 271144 3460
rect 252428 3420 271144 3448
rect 252428 3408 252434 3420
rect 271138 3408 271144 3420
rect 271196 3408 271202 3460
rect 413094 3448 413100 3460
rect 296686 3420 413100 3448
rect 30098 3340 30104 3392
rect 30156 3380 30162 3392
rect 40586 3380 40592 3392
rect 30156 3352 40592 3380
rect 30156 3340 30162 3352
rect 40586 3340 40592 3352
rect 40644 3340 40650 3392
rect 48958 3340 48964 3392
rect 49016 3380 49022 3392
rect 50338 3380 50344 3392
rect 49016 3352 50344 3380
rect 49016 3340 49022 3352
rect 50338 3340 50344 3352
rect 50396 3340 50402 3392
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 89254 3380 89260 3392
rect 84528 3352 89260 3380
rect 84528 3340 84534 3352
rect 89254 3340 89260 3352
rect 89312 3340 89318 3392
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 262950 3340 262956 3392
rect 263008 3380 263014 3392
rect 269850 3380 269856 3392
rect 263008 3352 269856 3380
rect 263008 3340 263014 3352
rect 269850 3340 269856 3352
rect 269908 3340 269914 3392
rect 292114 3340 292120 3392
rect 292172 3380 292178 3392
rect 296686 3380 296714 3420
rect 413094 3408 413100 3420
rect 413152 3408 413158 3460
rect 415486 3408 415492 3460
rect 415544 3448 415550 3460
rect 437566 3448 437572 3460
rect 415544 3420 437572 3448
rect 415544 3408 415550 3420
rect 437566 3408 437572 3420
rect 437624 3408 437630 3460
rect 450538 3408 450544 3460
rect 450596 3448 450602 3460
rect 452102 3448 452108 3460
rect 450596 3420 452108 3448
rect 450596 3408 450602 3420
rect 452102 3408 452108 3420
rect 452160 3408 452166 3460
rect 456886 3408 456892 3460
rect 456944 3448 456950 3460
rect 458082 3448 458088 3460
rect 456944 3420 458088 3448
rect 456944 3408 456950 3420
rect 458082 3408 458088 3420
rect 458140 3408 458146 3460
rect 569126 3448 569132 3460
rect 460906 3420 569132 3448
rect 292172 3352 296714 3380
rect 292172 3340 292178 3352
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332686 3340 332692 3392
rect 332744 3380 332750 3392
rect 333882 3380 333888 3392
rect 332744 3352 333888 3380
rect 332744 3340 332750 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 430850 3340 430856 3392
rect 430908 3380 430914 3392
rect 438026 3380 438032 3392
rect 430908 3352 438032 3380
rect 430908 3340 430914 3352
rect 438026 3340 438032 3352
rect 438084 3340 438090 3392
rect 445110 3340 445116 3392
rect 445168 3380 445174 3392
rect 460906 3380 460934 3420
rect 569126 3408 569132 3420
rect 569184 3408 569190 3460
rect 570598 3408 570604 3460
rect 570656 3448 570662 3460
rect 572714 3448 572720 3460
rect 570656 3420 572720 3448
rect 570656 3408 570662 3420
rect 572714 3408 572720 3420
rect 572772 3408 572778 3460
rect 445168 3352 460934 3380
rect 445168 3340 445174 3352
rect 57238 3272 57244 3324
rect 57296 3312 57302 3324
rect 58618 3312 58624 3324
rect 57296 3284 58624 3312
rect 57296 3272 57302 3284
rect 58618 3272 58624 3284
rect 58676 3272 58682 3324
rect 65518 3272 65524 3324
rect 65576 3312 65582 3324
rect 66898 3312 66904 3324
rect 65576 3284 66904 3312
rect 65576 3272 65582 3284
rect 66898 3272 66904 3284
rect 66956 3272 66962 3324
rect 259454 3272 259460 3324
rect 259512 3312 259518 3324
rect 264330 3312 264336 3324
rect 259512 3284 264336 3312
rect 259512 3272 259518 3284
rect 264330 3272 264336 3284
rect 264388 3272 264394 3324
rect 435542 3272 435548 3324
rect 435600 3312 435606 3324
rect 439314 3312 439320 3324
rect 435600 3284 439320 3312
rect 435600 3272 435606 3284
rect 439314 3272 439320 3284
rect 439372 3272 439378 3324
rect 6454 3204 6460 3256
rect 6512 3244 6518 3256
rect 7558 3244 7564 3256
rect 6512 3216 7564 3244
rect 6512 3204 6518 3216
rect 7558 3204 7564 3216
rect 7616 3204 7622 3256
rect 78582 3204 78588 3256
rect 78640 3244 78646 3256
rect 82170 3244 82176 3256
rect 78640 3216 82176 3244
rect 78640 3204 78646 3216
rect 82170 3204 82176 3216
rect 82228 3204 82234 3256
rect 478230 3204 478236 3256
rect 478288 3244 478294 3256
rect 479334 3244 479340 3256
rect 478288 3216 479340 3244
rect 478288 3204 478294 3216
rect 479334 3204 479340 3216
rect 479392 3204 479398 3256
rect 554038 3204 554044 3256
rect 554096 3244 554102 3256
rect 557350 3244 557356 3256
rect 554096 3216 557356 3244
rect 554096 3204 554102 3216
rect 557350 3204 557356 3216
rect 557408 3204 557414 3256
rect 293310 3136 293316 3188
rect 293368 3176 293374 3188
rect 296070 3176 296076 3188
rect 293368 3148 296076 3176
rect 293368 3136 293374 3148
rect 296070 3136 296076 3148
rect 296128 3136 296134 3188
rect 433242 3136 433248 3188
rect 433300 3176 433306 3188
rect 440418 3176 440424 3188
rect 433300 3148 440424 3176
rect 433300 3136 433306 3148
rect 440418 3136 440424 3148
rect 440476 3136 440482 3188
rect 485038 3136 485044 3188
rect 485096 3176 485102 3188
rect 487614 3176 487620 3188
rect 485096 3148 487620 3176
rect 485096 3136 485102 3148
rect 487614 3136 487620 3148
rect 487672 3136 487678 3188
rect 534718 3136 534724 3188
rect 534776 3176 534782 3188
rect 537202 3176 537208 3188
rect 534776 3148 537208 3176
rect 534776 3136 534782 3148
rect 537202 3136 537208 3148
rect 537260 3136 537266 3188
rect 560938 3136 560944 3188
rect 560996 3176 561002 3188
rect 563238 3176 563244 3188
rect 560996 3148 563244 3176
rect 560996 3136 561002 3148
rect 563238 3136 563244 3148
rect 563296 3136 563302 3188
rect 567838 3136 567844 3188
rect 567896 3176 567902 3188
rect 570322 3176 570328 3188
rect 567896 3148 570328 3176
rect 567896 3136 567902 3148
rect 570322 3136 570328 3148
rect 570380 3136 570386 3188
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 22738 3108 22744 3120
rect 19484 3080 22744 3108
rect 19484 3068 19490 3080
rect 22738 3068 22744 3080
rect 22796 3068 22802 3120
rect 273622 3068 273628 3120
rect 273680 3108 273686 3120
rect 278130 3108 278136 3120
rect 273680 3080 278136 3108
rect 273680 3068 273686 3080
rect 278130 3068 278136 3080
rect 278188 3068 278194 3120
rect 270034 3000 270040 3052
rect 270092 3040 270098 3052
rect 272518 3040 272524 3052
rect 270092 3012 272524 3040
rect 270092 3000 270098 3012
rect 272518 3000 272524 3012
rect 272576 3000 272582 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 472618 3000 472624 3052
rect 472676 3040 472682 3052
rect 474550 3040 474556 3052
rect 472676 3012 474556 3040
rect 472676 3000 472682 3012
rect 474550 3000 474556 3012
rect 474608 3000 474614 3052
rect 503070 3000 503076 3052
rect 503128 3040 503134 3052
rect 505370 3040 505376 3052
rect 503128 3012 505376 3040
rect 503128 3000 503134 3012
rect 505370 3000 505376 3012
rect 505428 3000 505434 3052
rect 538858 3000 538864 3052
rect 538916 3040 538922 3052
rect 540790 3040 540796 3052
rect 538916 3012 540796 3040
rect 538916 3000 538922 3012
rect 540790 3000 540796 3012
rect 540848 3000 540854 3052
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 565630 3040 565636 3052
rect 563756 3012 565636 3040
rect 563756 3000 563762 3012
rect 565630 3000 565636 3012
rect 565688 3000 565694 3052
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 14458 2972 14464 2984
rect 8812 2944 14464 2972
rect 8812 2932 8818 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 540238 2932 540244 2984
rect 540296 2972 540302 2984
rect 541986 2972 541992 2984
rect 540296 2944 541992 2972
rect 540296 2932 540302 2944
rect 541986 2932 541992 2944
rect 542044 2932 542050 2984
rect 552750 2932 552756 2984
rect 552808 2972 552814 2984
rect 554958 2972 554964 2984
rect 552808 2944 554964 2972
rect 552808 2932 552814 2944
rect 554958 2932 554964 2944
rect 555016 2932 555022 2984
rect 51350 2864 51356 2916
rect 51408 2904 51414 2916
rect 53098 2904 53104 2916
rect 51408 2876 53104 2904
rect 51408 2864 51414 2876
rect 53098 2864 53104 2876
rect 53156 2864 53162 2916
rect 73798 2864 73804 2916
rect 73856 2904 73862 2916
rect 75178 2904 75184 2916
rect 73856 2876 75184 2904
rect 73856 2864 73862 2876
rect 75178 2864 75184 2876
rect 75236 2864 75242 2916
rect 494790 2864 494796 2916
rect 494848 2904 494854 2916
rect 499390 2904 499396 2916
rect 494848 2876 499396 2904
rect 494848 2864 494854 2876
rect 499390 2864 499396 2876
rect 499448 2864 499454 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 348792 700544 348844 700596
rect 357624 700544 357676 700596
rect 332508 700476 332560 700528
rect 358912 700476 358964 700528
rect 300124 700408 300176 700460
rect 357532 700408 357584 700460
rect 283840 700340 283892 700392
rect 358820 700340 358872 700392
rect 105452 700272 105504 700324
rect 166264 700272 166316 700324
rect 217968 700272 218020 700324
rect 235172 700272 235224 700324
rect 267648 700272 267700 700324
rect 357440 700272 357492 700324
rect 371884 700272 371936 700324
rect 559656 700272 559708 700324
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 369124 696940 369176 696992
rect 580172 696940 580224 696992
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 3516 670692 3568 670744
rect 18604 670692 18656 670744
rect 360844 670692 360896 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 13084 656888 13136 656940
rect 373264 643084 373316 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 198004 632068 198056 632120
rect 377404 630640 377456 630692
rect 579988 630640 580040 630692
rect 378784 616836 378836 616888
rect 580172 616836 580224 616888
rect 3516 605820 3568 605872
rect 17224 605820 17276 605872
rect 363604 590656 363656 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 10324 579640 10376 579692
rect 367744 576852 367796 576904
rect 580172 576852 580224 576904
rect 359464 563048 359516 563100
rect 580172 563048 580224 563100
rect 3148 553664 3200 553716
rect 8944 553664 8996 553716
rect 500224 536800 500276 536852
rect 579896 536800 579948 536852
rect 2964 527144 3016 527196
rect 14464 527144 14516 527196
rect 2872 500964 2924 501016
rect 21364 500964 21416 501016
rect 482284 484372 482336 484424
rect 580172 484372 580224 484424
rect 217324 478864 217376 478916
rect 220084 478864 220136 478916
rect 217600 478252 217652 478304
rect 248420 478252 248472 478304
rect 309140 478252 309192 478304
rect 357624 478252 357676 478304
rect 218060 478184 218112 478236
rect 314752 478184 314804 478236
rect 71780 478116 71832 478168
rect 346492 478116 346544 478168
rect 217508 476756 217560 476808
rect 230480 476756 230532 476808
rect 238852 476756 238904 476808
rect 247040 476756 247092 476808
rect 237472 476688 237524 476740
rect 238760 476688 238812 476740
rect 233240 476620 233292 476672
rect 242900 476688 242952 476740
rect 291200 476688 291252 476740
rect 325792 476688 325844 476740
rect 233332 476552 233384 476604
rect 238852 476552 238904 476604
rect 236000 476416 236052 476468
rect 249800 476620 249852 476672
rect 251180 476620 251232 476672
rect 263600 476620 263652 476672
rect 278780 476620 278832 476672
rect 305000 476620 305052 476672
rect 248604 476552 248656 476604
rect 260840 476552 260892 476604
rect 280160 476552 280212 476604
rect 307760 476552 307812 476604
rect 242900 476484 242952 476536
rect 240140 476416 240192 476468
rect 231860 476280 231912 476332
rect 236000 476280 236052 476332
rect 236092 476280 236144 476332
rect 244280 476280 244332 476332
rect 238944 476212 238996 476264
rect 244372 476212 244424 476264
rect 245752 476484 245804 476536
rect 258264 476484 258316 476536
rect 259552 476484 259604 476536
rect 276020 476484 276072 476536
rect 281540 476484 281592 476536
rect 310520 476484 310572 476536
rect 255320 476416 255372 476468
rect 268016 476416 268068 476468
rect 282920 476416 282972 476468
rect 313280 476416 313332 476468
rect 247316 476280 247368 476332
rect 248512 476280 248564 476332
rect 252560 476348 252612 476400
rect 264980 476348 265032 476400
rect 284300 476348 284352 476400
rect 314660 476348 314712 476400
rect 255412 476280 255464 476332
rect 256792 476280 256844 476332
rect 270500 476280 270552 476332
rect 285680 476280 285732 476332
rect 317420 476280 317472 476332
rect 252744 476212 252796 476264
rect 258172 476212 258224 476264
rect 273260 476212 273312 476264
rect 288440 476212 288492 476264
rect 320180 476212 320232 476264
rect 234620 476144 234672 476196
rect 237380 476144 237432 476196
rect 241520 476144 241572 476196
rect 245660 476144 245712 476196
rect 253848 476144 253900 476196
rect 256700 476144 256752 476196
rect 260932 476144 260984 476196
rect 277952 476144 278004 476196
rect 289820 476144 289872 476196
rect 322940 476144 322992 476196
rect 234712 476076 234764 476128
rect 236000 476076 236052 476128
rect 242808 476076 242860 476128
rect 244280 476076 244332 476128
rect 245844 476076 245896 476128
rect 247040 476076 247092 476128
rect 252468 476076 252520 476128
rect 253940 476076 253992 476128
rect 258080 476076 258132 476128
rect 262220 476076 262272 476128
rect 277584 476076 277636 476128
rect 302240 476076 302292 476128
rect 219072 475328 219124 475380
rect 238852 475328 238904 475380
rect 267556 475328 267608 475380
rect 274640 475328 274692 475380
rect 3332 474716 3384 474768
rect 331220 474716 331272 474768
rect 219164 474036 219216 474088
rect 241612 474036 241664 474088
rect 274456 474036 274508 474088
rect 284392 474036 284444 474088
rect 298100 474036 298152 474088
rect 377404 474036 377456 474088
rect 198004 473968 198056 474020
rect 324320 473968 324372 474020
rect 217784 472676 217836 472728
rect 251272 472676 251324 472728
rect 14464 472608 14516 472660
rect 328460 472608 328512 472660
rect 217876 471316 217928 471368
rect 254032 471316 254084 471368
rect 6920 471248 6972 471300
rect 347872 471248 347924 471300
rect 300860 469888 300912 469940
rect 580264 469888 580316 469940
rect 10324 469820 10376 469872
rect 327080 469820 327132 469872
rect 166264 468460 166316 468512
rect 317420 468460 317472 468512
rect 320180 468460 320232 468512
rect 500224 468460 500276 468512
rect 295340 467168 295392 467220
rect 367744 467168 367796 467220
rect 4804 467100 4856 467152
rect 321560 467100 321612 467152
rect 276020 465740 276072 465792
rect 300952 465740 301004 465792
rect 169760 465672 169812 465724
rect 314752 465672 314804 465724
rect 318800 465672 318852 465724
rect 482284 465672 482336 465724
rect 273260 464380 273312 464432
rect 298192 464380 298244 464432
rect 307760 464380 307812 464432
rect 364340 464380 364392 464432
rect 17224 464312 17276 464364
rect 350540 464312 350592 464364
rect 266452 462952 266504 463004
rect 285772 462952 285824 463004
rect 3332 462340 3384 462392
rect 332600 462340 332652 462392
rect 275928 461660 275980 461712
rect 285772 461660 285824 461712
rect 219256 461592 219308 461644
rect 244372 461592 244424 461644
rect 263692 461592 263744 461644
rect 280252 461592 280304 461644
rect 325700 461592 325752 461644
rect 373264 461592 373316 461644
rect 271880 460232 271932 460284
rect 295432 460232 295484 460284
rect 322940 460232 322992 460284
rect 363604 460232 363656 460284
rect 13084 460164 13136 460216
rect 350632 460164 350684 460216
rect 269488 458872 269540 458924
rect 289912 458872 289964 458924
rect 306380 458872 306432 458924
rect 428464 458872 428516 458924
rect 8944 458804 8996 458856
rect 351920 458804 351972 458856
rect 268016 457512 268068 457564
rect 287060 457512 287112 457564
rect 303712 457512 303764 457564
rect 494060 457512 494112 457564
rect 21364 457444 21416 457496
rect 352472 457444 352524 457496
rect 265072 456084 265124 456136
rect 283012 456084 283064 456136
rect 301320 456084 301372 456136
rect 371884 456084 371936 456136
rect 18604 456016 18656 456068
rect 323768 456016 323820 456068
rect 269028 455336 269080 455388
rect 276480 455336 276532 455388
rect 274548 454724 274600 454776
rect 283012 454724 283064 454776
rect 219348 454656 219400 454708
rect 247132 454656 247184 454708
rect 280068 454656 280120 454708
rect 290464 454656 290516 454708
rect 298928 454656 298980 454708
rect 360844 454656 360896 454708
rect 267648 453364 267700 453416
rect 273352 453364 273404 453416
rect 277308 453364 277360 453416
rect 287336 453364 287388 453416
rect 270960 453296 271012 453348
rect 292580 453296 292632 453348
rect 296720 453296 296772 453348
rect 378784 453296 378836 453348
rect 271788 452752 271840 452804
rect 279608 452752 279660 452804
rect 266268 451936 266320 451988
rect 271972 451936 272024 451988
rect 273168 451936 273220 451988
rect 281724 451936 281776 451988
rect 217692 451868 217744 451920
rect 231952 451868 232004 451920
rect 270408 451868 270460 451920
rect 277492 451868 277544 451920
rect 278688 451868 278740 451920
rect 288808 451868 288860 451920
rect 294328 451868 294380 451920
rect 359464 451868 359516 451920
rect 328092 450644 328144 450696
rect 369124 450644 369176 450696
rect 3516 450576 3568 450628
rect 328828 450576 328880 450628
rect 3608 450508 3660 450560
rect 331220 450508 331272 450560
rect 307944 449556 307996 449608
rect 412640 449556 412692 449608
rect 153200 449488 153252 449540
rect 317236 449488 317288 449540
rect 305552 449420 305604 449472
rect 477500 449420 477552 449472
rect 88340 449352 88392 449404
rect 319536 449352 319588 449404
rect 303252 449284 303304 449336
rect 542360 449284 542412 449336
rect 23480 449216 23532 449268
rect 321836 449216 321888 449268
rect 3424 449148 3476 449200
rect 326528 449148 326580 449200
rect 335084 448128 335136 448180
rect 397460 448128 397512 448180
rect 332784 448060 332836 448112
rect 462320 448060 462372 448112
rect 201500 447992 201552 448044
rect 342076 447992 342128 448044
rect 136640 447924 136692 447976
rect 344376 447924 344428 447976
rect 40040 447856 40092 447908
rect 320364 447856 320416 447908
rect 330392 447856 330444 447908
rect 527180 447856 527232 447908
rect 2872 447788 2924 447840
rect 353668 447788 353720 447840
rect 231860 447040 231912 447092
rect 232412 447040 232464 447092
rect 236000 447040 236052 447092
rect 237012 447040 237064 447092
rect 241520 447040 241572 447092
rect 242348 447040 242400 447092
rect 245752 447040 245804 447092
rect 246396 447040 246448 447092
rect 248420 447040 248472 447092
rect 249340 447040 249392 447092
rect 252560 447040 252612 447092
rect 253204 447040 253256 447092
rect 255964 447040 256016 447092
rect 258264 447040 258316 447092
rect 258724 447040 258776 447092
rect 261116 447040 261168 447092
rect 262864 447040 262916 447092
rect 267556 447040 267608 447092
rect 271880 447040 271932 447092
rect 272708 447040 272760 447092
rect 273260 447040 273312 447092
rect 274180 447040 274232 447092
rect 277492 447040 277544 447092
rect 278044 447040 278096 447092
rect 281540 447040 281592 447092
rect 281908 447040 281960 447092
rect 282920 447040 282972 447092
rect 283564 447040 283616 447092
rect 284300 447040 284352 447092
rect 285036 447040 285088 447092
rect 285680 447040 285732 447092
rect 286692 447040 286744 447092
rect 350540 447040 350592 447092
rect 351092 447040 351144 447092
rect 256608 446972 256660 447024
rect 259828 446972 259880 447024
rect 260748 446972 260800 447024
rect 264520 446972 264572 447024
rect 264244 446904 264296 446956
rect 269120 446904 269172 446956
rect 57244 446768 57296 446820
rect 349804 446768 349856 446820
rect 339684 446700 339736 446752
rect 357440 446700 357492 446752
rect 217968 446632 218020 446684
rect 313372 446632 313424 446684
rect 337384 446632 337436 446684
rect 358912 446632 358964 446684
rect 312544 446564 312596 446616
rect 358820 446564 358872 446616
rect 261484 446496 261536 446548
rect 265992 446496 266044 446548
rect 310980 446496 311032 446548
rect 357532 446496 357584 446548
rect 220084 446428 220136 446480
rect 230388 446428 230440 446480
rect 265624 446428 265676 446480
rect 270684 446428 270736 446480
rect 307116 446428 307168 446480
rect 364984 446428 365036 446480
rect 311808 446360 311860 446412
rect 362224 446360 362276 446412
rect 304816 446292 304868 446344
rect 363604 446292 363656 446344
rect 293132 446224 293184 446276
rect 362316 446224 362368 446276
rect 292396 446156 292448 446208
rect 373264 446156 373316 446208
rect 244372 446088 244424 446140
rect 345112 446088 345164 446140
rect 229836 446020 229888 446072
rect 338212 446020 338264 446072
rect 228364 445952 228416 446004
rect 347504 445952 347556 446004
rect 229744 445884 229796 445936
rect 359924 445884 359976 445936
rect 293960 445816 294012 445868
rect 458824 445816 458876 445868
rect 302516 445748 302568 445800
rect 311164 445748 311216 445800
rect 316408 445748 316460 445800
rect 333980 445748 334032 445800
rect 253940 445408 253992 445460
rect 254860 445408 254912 445460
rect 228548 445204 228600 445256
rect 336648 445204 336700 445256
rect 225696 445136 225748 445188
rect 338948 445136 339000 445188
rect 333980 445068 334032 445120
rect 580356 445068 580408 445120
rect 311164 445000 311216 445052
rect 580264 445000 580316 445052
rect 224224 444932 224276 444984
rect 341248 444932 341300 444984
rect 228456 444864 228508 444916
rect 355968 444864 356020 444916
rect 300124 444796 300176 444848
rect 460204 444796 460256 444848
rect 295524 444728 295576 444780
rect 494704 444728 494756 444780
rect 86224 444660 86276 444712
rect 343640 444660 343692 444712
rect 84844 444592 84896 444644
rect 345940 444592 345992 444644
rect 82084 444524 82136 444576
rect 348240 444524 348292 444576
rect 80704 444456 80756 444508
rect 358360 444456 358412 444508
rect 7564 444388 7616 444440
rect 334256 444388 334308 444440
rect 309508 443708 309560 443760
rect 3516 443640 3568 443692
rect 244372 443640 244424 443692
rect 314384 443640 314436 443692
rect 369124 443640 369176 443692
rect 367744 443572 367796 443624
rect 226984 443504 227036 443556
rect 335544 443504 335596 443556
rect 225604 443436 225656 443488
rect 340236 443436 340288 443488
rect 220084 443368 220136 443420
rect 342444 443368 342496 443420
rect 228640 443300 228692 443352
rect 354220 443300 354272 443352
rect 221464 443232 221516 443284
rect 354956 443232 355008 443284
rect 298008 443164 298060 443216
rect 446404 443164 446456 443216
rect 98644 443096 98696 443148
rect 356428 443096 356480 443148
rect 95976 443028 96028 443080
rect 357440 443028 357492 443080
rect 358820 443028 358872 443080
rect 79324 442960 79376 443012
rect 3608 442212 3660 442264
rect 229836 442212 229888 442264
rect 362316 439492 362368 439544
rect 581000 439492 581052 439544
rect 458824 438132 458876 438184
rect 582380 438132 582432 438184
rect 3424 423580 3476 423632
rect 7564 423580 7616 423632
rect 2964 411204 3016 411256
rect 226984 411204 227036 411256
rect 3424 410524 3476 410576
rect 229744 410524 229796 410576
rect 3332 398760 3384 398812
rect 228640 398760 228692 398812
rect 369124 379448 369176 379500
rect 580172 379448 580224 379500
rect 3056 372512 3108 372564
rect 228548 372512 228600 372564
rect 3332 346332 3384 346384
rect 221464 346332 221516 346384
rect 362224 325592 362276 325644
rect 579896 325592 579948 325644
rect 3332 320084 3384 320136
rect 225696 320084 225748 320136
rect 261024 310496 261076 310548
rect 261208 310496 261260 310548
rect 266544 310496 266596 310548
rect 266728 310496 266780 310548
rect 291476 310496 291528 310548
rect 291660 310496 291712 310548
rect 292764 310496 292816 310548
rect 292948 310496 293000 310548
rect 300860 310496 300912 310548
rect 301228 310496 301280 310548
rect 310612 310496 310664 310548
rect 310796 310496 310848 310548
rect 327356 310496 327408 310548
rect 327540 310496 327592 310548
rect 353484 310496 353536 310548
rect 353668 310496 353720 310548
rect 44824 309748 44876 309800
rect 361120 309748 361172 309800
rect 229652 309068 229704 309120
rect 236552 309068 236604 309120
rect 284116 309068 284168 309120
rect 338580 309068 338632 309120
rect 342168 309068 342220 309120
rect 342904 309068 342956 309120
rect 95884 308932 95936 308984
rect 237196 309000 237248 309052
rect 290280 309000 290332 309052
rect 293500 309000 293552 309052
rect 296260 309000 296312 309052
rect 352932 309000 352984 309052
rect 229744 308932 229796 308984
rect 235908 308932 235960 308984
rect 97264 308864 97316 308916
rect 247684 308932 247736 308984
rect 286416 308932 286468 308984
rect 350908 308932 350960 308984
rect 355048 308932 355100 308984
rect 282828 308864 282880 308916
rect 348148 308864 348200 308916
rect 71044 308796 71096 308848
rect 234620 308796 234672 308848
rect 242256 308796 242308 308848
rect 260932 308796 260984 308848
rect 283932 308796 283984 308848
rect 352012 308796 352064 308848
rect 64144 308728 64196 308780
rect 232872 308728 232924 308780
rect 235816 308728 235868 308780
rect 243728 308728 243780 308780
rect 275560 308728 275612 308780
rect 279884 308728 279936 308780
rect 285588 308728 285640 308780
rect 354036 308728 354088 308780
rect 46204 308660 46256 308712
rect 229652 308660 229704 308712
rect 257344 308660 257396 308712
rect 277032 308660 277084 308712
rect 287704 308660 287756 308712
rect 348792 308660 348844 308712
rect 354404 308660 354456 308712
rect 355692 308728 355744 308780
rect 31760 308592 31812 308644
rect 229744 308592 229796 308644
rect 243728 308592 243780 308644
rect 251180 308592 251232 308644
rect 253572 308592 253624 308644
rect 254400 308592 254452 308644
rect 279884 308592 279936 308644
rect 349436 308592 349488 308644
rect 356244 308592 356296 308644
rect 356428 308592 356480 308644
rect 359004 308592 359056 308644
rect 359280 308592 359332 308644
rect 438032 308728 438084 308780
rect 436836 308660 436888 308712
rect 439504 308592 439556 308644
rect 39304 308524 39356 308576
rect 232044 308524 232096 308576
rect 249064 308524 249116 308576
rect 347688 308524 347740 308576
rect 353760 308524 353812 308576
rect 439596 308524 439648 308576
rect 27620 308456 27672 308508
rect 235264 308456 235316 308508
rect 236828 308456 236880 308508
rect 246396 308456 246448 308508
rect 247684 308456 247736 308508
rect 348976 308456 349028 308508
rect 353116 308456 353168 308508
rect 438124 308456 438176 308508
rect 23480 308388 23532 308440
rect 234436 308388 234488 308440
rect 238024 308388 238076 308440
rect 282644 308320 282696 308372
rect 283656 308320 283708 308372
rect 340880 308388 340932 308440
rect 341892 308388 341944 308440
rect 342536 308388 342588 308440
rect 343180 308388 343232 308440
rect 343640 308388 343692 308440
rect 343916 308388 343968 308440
rect 345204 308388 345256 308440
rect 345940 308388 345992 308440
rect 346584 308388 346636 308440
rect 346860 308388 346912 308440
rect 349344 308388 349396 308440
rect 350080 308388 350132 308440
rect 352472 308388 352524 308440
rect 440516 308388 440568 308440
rect 250444 308184 250496 308236
rect 252652 308184 252704 308236
rect 281448 308184 281500 308236
rect 283748 308184 283800 308236
rect 247592 308116 247644 308168
rect 252284 308116 252336 308168
rect 243636 308048 243688 308100
rect 250076 308048 250128 308100
rect 252652 308048 252704 308100
rect 253296 308048 253348 308100
rect 283748 308048 283800 308100
rect 337476 308252 337528 308304
rect 341156 308252 341208 308304
rect 341800 308252 341852 308304
rect 342628 308252 342680 308304
rect 343548 308252 343600 308304
rect 320180 308184 320232 308236
rect 320732 308184 320784 308236
rect 342352 308184 342404 308236
rect 343088 308184 343140 308236
rect 345112 308320 345164 308372
rect 345572 308320 345624 308372
rect 346676 308320 346728 308372
rect 347228 308320 347280 308372
rect 354680 308320 354732 308372
rect 354864 308320 354916 308372
rect 356152 308320 356204 308372
rect 356796 308320 356848 308372
rect 357532 308320 357584 308372
rect 358084 308320 358136 308372
rect 345296 308252 345348 308304
rect 345480 308252 345532 308304
rect 356060 308252 356112 308304
rect 357256 308252 357308 308304
rect 357716 308252 357768 308304
rect 358176 308252 358228 308304
rect 359188 308252 359240 308304
rect 359832 308252 359884 308304
rect 360200 308252 360252 308304
rect 360476 308252 360528 308304
rect 350264 308184 350316 308236
rect 357624 308184 357676 308236
rect 358544 308184 358596 308236
rect 359096 308184 359148 308236
rect 359924 308184 359976 308236
rect 284392 308048 284444 308100
rect 293224 308048 293276 308100
rect 246396 307980 246448 308032
rect 250260 307980 250312 308032
rect 283564 307980 283616 308032
rect 285220 307980 285272 308032
rect 246856 307912 246908 307964
rect 249892 307912 249944 307964
rect 261208 307912 261260 307964
rect 261668 307912 261720 307964
rect 274088 307912 274140 307964
rect 279424 307912 279476 307964
rect 279792 307912 279844 307964
rect 287704 307912 287756 307964
rect 291016 307912 291068 307964
rect 337660 308116 337712 308168
rect 345296 308116 345348 308168
rect 346124 308116 346176 308168
rect 350816 308116 350868 308168
rect 351460 308116 351512 308168
rect 354772 308116 354824 308168
rect 355508 308116 355560 308168
rect 358820 308116 358872 308168
rect 359464 308116 359516 308168
rect 350632 308048 350684 308100
rect 351368 308048 351420 308100
rect 359280 308048 359332 308100
rect 240876 307844 240928 307896
rect 229744 307776 229796 307828
rect 230940 307776 230992 307828
rect 236736 307776 236788 307828
rect 238116 307776 238168 307828
rect 239772 307776 239824 307828
rect 241152 307776 241204 307828
rect 242164 307776 242216 307828
rect 242900 307776 242952 307828
rect 246304 307844 246356 307896
rect 248972 307844 249024 307896
rect 253388 307844 253440 307896
rect 259644 307844 259696 307896
rect 260104 307844 260156 307896
rect 262864 307844 262916 307896
rect 268476 307844 268528 307896
rect 275744 307844 275796 307896
rect 278872 307844 278924 307896
rect 281356 307844 281408 307896
rect 284668 307844 284720 307896
rect 286324 307844 286376 307896
rect 293960 307844 294012 307896
rect 295800 307844 295852 307896
rect 317512 307844 317564 307896
rect 320824 307844 320876 307896
rect 334256 307844 334308 307896
rect 334808 307844 334860 307896
rect 359372 307844 359424 307896
rect 247684 307776 247736 307828
rect 247776 307776 247828 307828
rect 248512 307776 248564 307828
rect 253296 307776 253348 307828
rect 253572 307776 253624 307828
rect 254952 307776 255004 307828
rect 255688 307776 255740 307828
rect 256240 307776 256292 307828
rect 258356 307776 258408 307828
rect 261668 307776 261720 307828
rect 262220 307776 262272 307828
rect 265624 307776 265676 307828
rect 266820 307776 266872 307828
rect 269764 307776 269816 307828
rect 272064 307776 272116 307828
rect 278044 307776 278096 307828
rect 278964 307776 279016 307828
rect 279700 307776 279752 307828
rect 281172 307776 281224 307828
rect 284024 307776 284076 307828
rect 284944 307776 284996 307828
rect 286784 307776 286836 307828
rect 289084 307776 289136 307828
rect 292672 307776 292724 307828
rect 294512 307776 294564 307828
rect 295248 307776 295300 307828
rect 296076 307776 296128 307828
rect 314844 307776 314896 307828
rect 318064 307776 318116 307828
rect 343640 307232 343692 307284
rect 344652 307232 344704 307284
rect 68284 307164 68336 307216
rect 241796 307164 241848 307216
rect 334624 307164 334676 307216
rect 445024 307164 445076 307216
rect 57980 307096 58032 307148
rect 240692 307096 240744 307148
rect 318340 307096 318392 307148
rect 462964 307096 463016 307148
rect 25504 307028 25556 307080
rect 230112 307028 230164 307080
rect 238024 307028 238076 307080
rect 252928 307028 252980 307080
rect 264244 307028 264296 307080
rect 274640 307028 274692 307080
rect 322204 307028 322256 307080
rect 500224 307028 500276 307080
rect 257068 306960 257120 307012
rect 268108 306960 268160 307012
rect 287244 306960 287296 307012
rect 257160 306756 257212 306808
rect 268200 306756 268252 306808
rect 287336 306756 287388 306808
rect 233516 306688 233568 306740
rect 259828 306688 259880 306740
rect 233516 306484 233568 306536
rect 238760 306484 238812 306536
rect 239128 306484 239180 306536
rect 245660 306484 245712 306536
rect 245936 306484 245988 306536
rect 320272 306620 320324 306672
rect 321100 306620 321152 306672
rect 303804 306552 303856 306604
rect 304356 306552 304408 306604
rect 325792 306552 325844 306604
rect 326804 306552 326856 306604
rect 350724 306552 350776 306604
rect 351828 306552 351880 306604
rect 287152 306484 287204 306536
rect 287428 306484 287480 306536
rect 292672 306484 292724 306536
rect 293776 306484 293828 306536
rect 294052 306484 294104 306536
rect 295064 306484 295116 306536
rect 295432 306484 295484 306536
rect 296168 306484 296220 306536
rect 299572 306484 299624 306536
rect 300124 306484 300176 306536
rect 302424 306484 302476 306536
rect 303344 306484 303396 306536
rect 313740 306484 313792 306536
rect 313924 306484 313976 306536
rect 316132 306484 316184 306536
rect 317236 306484 317288 306536
rect 320272 306484 320324 306536
rect 321008 306484 321060 306536
rect 325884 306484 325936 306536
rect 326252 306484 326304 306536
rect 327172 306484 327224 306536
rect 328184 306484 328236 306536
rect 331220 306484 331272 306536
rect 331772 306484 331824 306536
rect 333980 306484 334032 306536
rect 334532 306484 334584 306536
rect 234712 306416 234764 306468
rect 235356 306416 235408 306468
rect 232044 306348 232096 306400
rect 232964 306348 233016 306400
rect 3332 306280 3384 306332
rect 225604 306280 225656 306332
rect 229192 306280 229244 306332
rect 230296 306280 230348 306332
rect 231952 306280 232004 306332
rect 232504 306280 232556 306332
rect 236184 306280 236236 306332
rect 237012 306280 237064 306332
rect 239404 306416 239456 306468
rect 245844 306416 245896 306468
rect 246580 306416 246632 306468
rect 259828 306416 259880 306468
rect 272064 306416 272116 306468
rect 272892 306416 272944 306468
rect 273444 306416 273496 306468
rect 273628 306416 273680 306468
rect 281632 306416 281684 306468
rect 282184 306416 282236 306468
rect 285680 306416 285732 306468
rect 286600 306416 286652 306468
rect 287060 306416 287112 306468
rect 287612 306416 287664 306468
rect 288532 306416 288584 306468
rect 288808 306416 288860 306468
rect 292580 306416 292632 306468
rect 293316 306416 293368 306468
rect 293960 306416 294012 306468
rect 294420 306416 294472 306468
rect 295616 306416 295668 306468
rect 296352 306416 296404 306468
rect 299480 306416 299532 306468
rect 300032 306416 300084 306468
rect 302240 306416 302292 306468
rect 302700 306416 302752 306468
rect 306472 306416 306524 306468
rect 306748 306416 306800 306468
rect 312268 306416 312320 306468
rect 312636 306416 312688 306468
rect 313280 306416 313332 306468
rect 314200 306416 314252 306468
rect 316040 306416 316092 306468
rect 316776 306416 316828 306468
rect 322940 306416 322992 306468
rect 323492 306416 323544 306468
rect 325700 306416 325752 306468
rect 326160 306416 326212 306468
rect 327080 306416 327132 306468
rect 327908 306416 327960 306468
rect 329840 306416 329892 306468
rect 330668 306416 330720 306468
rect 241796 306348 241848 306400
rect 242532 306348 242584 306400
rect 247408 306348 247460 306400
rect 248328 306348 248380 306400
rect 248512 306348 248564 306400
rect 249248 306348 249300 306400
rect 259552 306348 259604 306400
rect 260564 306348 260616 306400
rect 262404 306348 262456 306400
rect 262956 306348 263008 306400
rect 266820 306348 266872 306400
rect 267464 306348 267516 306400
rect 267740 306348 267792 306400
rect 268384 306348 268436 306400
rect 269396 306348 269448 306400
rect 270040 306348 270092 306400
rect 272156 306348 272208 306400
rect 272524 306348 272576 306400
rect 285772 306348 285824 306400
rect 286140 306348 286192 306400
rect 287428 306348 287480 306400
rect 288164 306348 288216 306400
rect 288440 306348 288492 306400
rect 289268 306348 289320 306400
rect 289820 306348 289872 306400
rect 290096 306348 290148 306400
rect 291200 306348 291252 306400
rect 291568 306348 291620 306400
rect 291660 306348 291712 306400
rect 292212 306348 292264 306400
rect 292856 306348 292908 306400
rect 293408 306348 293460 306400
rect 294144 306348 294196 306400
rect 294604 306348 294656 306400
rect 295524 306348 295576 306400
rect 295984 306348 296036 306400
rect 296720 306348 296772 306400
rect 297456 306348 297508 306400
rect 298100 306348 298152 306400
rect 298560 306348 298612 306400
rect 299756 306348 299808 306400
rect 300584 306348 300636 306400
rect 301228 306348 301280 306400
rect 301780 306348 301832 306400
rect 302516 306348 302568 306400
rect 302884 306348 302936 306400
rect 303712 306348 303764 306400
rect 304632 306348 304684 306400
rect 306564 306348 306616 306400
rect 307208 306348 307260 306400
rect 307760 306348 307812 306400
rect 308404 306348 308456 306400
rect 309140 306348 309192 306400
rect 310060 306348 310112 306400
rect 310704 306348 310756 306400
rect 311808 306348 311860 306400
rect 313464 306348 313516 306400
rect 314384 306348 314436 306400
rect 314844 306348 314896 306400
rect 315304 306348 315356 306400
rect 316224 306348 316276 306400
rect 316868 306348 316920 306400
rect 317420 306348 317472 306400
rect 317972 306348 318024 306400
rect 318892 306348 318944 306400
rect 319812 306348 319864 306400
rect 320456 306348 320508 306400
rect 321376 306348 321428 306400
rect 324320 306348 324372 306400
rect 325056 306348 325108 306400
rect 325884 306348 325936 306400
rect 326436 306348 326488 306400
rect 327448 306348 327500 306400
rect 328092 306348 328144 306400
rect 328460 306348 328512 306400
rect 329196 306348 329248 306400
rect 241704 306280 241756 306332
rect 242440 306280 242492 306332
rect 247316 306280 247368 306332
rect 247868 306280 247920 306332
rect 248696 306280 248748 306332
rect 249156 306280 249208 306332
rect 249892 306280 249944 306332
rect 250720 306280 250772 306332
rect 252744 306280 252796 306332
rect 253756 306280 253808 306332
rect 254216 306280 254268 306332
rect 255044 306280 255096 306332
rect 255780 306280 255832 306332
rect 256332 306280 256384 306332
rect 256884 306280 256936 306332
rect 257436 306280 257488 306332
rect 258172 306280 258224 306332
rect 259184 306280 259236 306332
rect 259736 306280 259788 306332
rect 260472 306280 260524 306332
rect 262588 306280 262640 306332
rect 263508 306280 263560 306332
rect 263692 306280 263744 306332
rect 263968 306280 264020 306332
rect 265348 306280 265400 306332
rect 265992 306280 266044 306332
rect 266636 306280 266688 306332
rect 267004 306280 267056 306332
rect 268016 306280 268068 306332
rect 268844 306280 268896 306332
rect 269304 306280 269356 306332
rect 269856 306280 269908 306332
rect 271972 306280 272024 306332
rect 272432 306280 272484 306332
rect 273260 306280 273312 306332
rect 274180 306280 274232 306332
rect 274732 306280 274784 306332
rect 274916 306280 274968 306332
rect 277400 306280 277452 306332
rect 278504 306280 278556 306332
rect 280436 306280 280488 306332
rect 280896 306280 280948 306332
rect 280988 306280 281040 306332
rect 331956 306416 332008 306468
rect 332692 306416 332744 306468
rect 333060 306416 333112 306468
rect 333980 306348 334032 306400
rect 335084 306348 335136 306400
rect 335636 306348 335688 306400
rect 336556 306348 336608 306400
rect 331312 306280 331364 306332
rect 332324 306280 332376 306332
rect 332600 306280 332652 306332
rect 333612 306280 333664 306332
rect 334072 306280 334124 306332
rect 334716 306280 334768 306332
rect 335728 306280 335780 306332
rect 336004 306280 336056 306332
rect 336924 306280 336976 306332
rect 337108 306280 337160 306332
rect 338212 306280 338264 306332
rect 339408 306280 339460 306332
rect 339592 306280 339644 306332
rect 340696 306280 340748 306332
rect 230940 306212 230992 306264
rect 231584 306212 231636 306264
rect 237472 306212 237524 306264
rect 237932 306212 237984 306264
rect 238852 306212 238904 306264
rect 239036 306212 239088 306264
rect 239680 306212 239732 306264
rect 240416 306212 240468 306264
rect 241336 306212 241388 306264
rect 243176 306212 243228 306264
rect 244188 306212 244240 306264
rect 244740 306212 244792 306264
rect 245476 306212 245528 306264
rect 246028 306212 246080 306264
rect 246764 306212 246816 306264
rect 247500 306212 247552 306264
rect 247960 306212 248012 306264
rect 250076 306212 250128 306264
rect 250904 306212 250956 306264
rect 262312 306212 262364 306264
rect 263324 306212 263376 306264
rect 265256 306212 265308 306264
rect 265716 306212 265768 306264
rect 266544 306212 266596 306264
rect 267648 306212 267700 306264
rect 268108 306212 268160 306264
rect 268752 306212 268804 306264
rect 269212 306212 269264 306264
rect 270132 306212 270184 306264
rect 270684 306212 270736 306264
rect 271052 306212 271104 306264
rect 273352 306212 273404 306264
rect 273720 306212 273772 306264
rect 277584 306212 277636 306264
rect 278320 306212 278372 306264
rect 237748 306144 237800 306196
rect 238392 306144 238444 306196
rect 238760 306144 238812 306196
rect 240048 306144 240100 306196
rect 257068 306144 257120 306196
rect 257528 306144 257580 306196
rect 258356 306144 258408 306196
rect 258816 306144 258868 306196
rect 259460 306144 259512 306196
rect 260012 306144 260064 306196
rect 270868 306144 270920 306196
rect 274916 306144 274968 306196
rect 275928 306144 275980 306196
rect 276940 306144 276992 306196
rect 340972 306212 341024 306264
rect 237564 306076 237616 306128
rect 238300 306076 238352 306128
rect 255504 306076 255556 306128
rect 255964 306076 256016 306128
rect 256792 306076 256844 306128
rect 257896 306076 257948 306128
rect 263968 306076 264020 306128
rect 264704 306076 264756 306128
rect 255412 306008 255464 306060
rect 256424 306008 256476 306060
rect 230848 305940 230900 305992
rect 231124 305940 231176 305992
rect 263784 305940 263836 305992
rect 264428 305940 264480 305992
rect 270592 305940 270644 305992
rect 277032 306076 277084 306128
rect 342260 306144 342312 306196
rect 277124 306008 277176 306060
rect 280988 306076 281040 306128
rect 281724 306076 281776 306128
rect 282460 306076 282512 306128
rect 282736 306076 282788 306128
rect 350632 306076 350684 306128
rect 282644 306008 282696 306060
rect 354864 306008 354916 306060
rect 281080 305940 281132 305992
rect 354220 305940 354272 305992
rect 270684 305872 270736 305924
rect 271604 305872 271656 305924
rect 280988 305872 281040 305924
rect 354680 305872 354732 305924
rect 270500 305804 270552 305856
rect 271788 305804 271840 305856
rect 280896 305804 280948 305856
rect 354772 305804 354824 305856
rect 280804 305736 280856 305788
rect 356152 305736 356204 305788
rect 75920 305668 75972 305720
rect 244004 305668 244056 305720
rect 277308 305668 277360 305720
rect 353668 305668 353720 305720
rect 72424 305600 72476 305652
rect 242992 305600 243044 305652
rect 278320 305600 278372 305652
rect 357440 305600 357492 305652
rect 283012 305532 283064 305584
rect 284208 305532 284260 305584
rect 284392 305532 284444 305584
rect 285128 305532 285180 305584
rect 287244 305532 287296 305584
rect 287888 305532 287940 305584
rect 288624 305532 288676 305584
rect 289176 305532 289228 305584
rect 290004 305532 290056 305584
rect 290464 305532 290516 305584
rect 291200 305532 291252 305584
rect 292028 305532 292080 305584
rect 284484 305464 284536 305516
rect 285036 305464 285088 305516
rect 287060 305464 287112 305516
rect 288072 305464 288124 305516
rect 288808 305464 288860 305516
rect 289636 305464 289688 305516
rect 289820 305464 289872 305516
rect 290556 305464 290608 305516
rect 283932 305396 283984 305448
rect 284208 305396 284260 305448
rect 289544 305396 289596 305448
rect 332508 305532 332560 305584
rect 332876 305532 332928 305584
rect 333336 305532 333388 305584
rect 334256 305532 334308 305584
rect 335268 305532 335320 305584
rect 335544 305532 335596 305584
rect 336372 305532 336424 305584
rect 339684 305532 339736 305584
rect 340144 305532 340196 305584
rect 294236 305464 294288 305516
rect 294696 305464 294748 305516
rect 295800 305464 295852 305516
rect 295984 305464 296036 305516
rect 299848 305464 299900 305516
rect 300492 305464 300544 305516
rect 300952 305464 301004 305516
rect 301596 305464 301648 305516
rect 301044 305396 301096 305448
rect 301872 305396 301924 305448
rect 236644 305328 236696 305380
rect 236828 305328 236880 305380
rect 295064 305260 295116 305312
rect 340880 305464 340932 305516
rect 260932 305192 260984 305244
rect 262036 305192 262088 305244
rect 298008 305192 298060 305244
rect 303804 305328 303856 305380
rect 304816 305328 304868 305380
rect 305276 305328 305328 305380
rect 306012 305328 306064 305380
rect 306380 305328 306432 305380
rect 306840 305328 306892 305380
rect 308036 305328 308088 305380
rect 308772 305328 308824 305380
rect 309324 305328 309376 305380
rect 309692 305328 309744 305380
rect 310520 305328 310572 305380
rect 310888 305328 310940 305380
rect 311992 305328 312044 305380
rect 313096 305328 313148 305380
rect 313556 305328 313608 305380
rect 313832 305328 313884 305380
rect 314936 305328 314988 305380
rect 315580 305328 315632 305380
rect 317696 305328 317748 305380
rect 318524 305328 318576 305380
rect 318800 305328 318852 305380
rect 319168 305328 319220 305380
rect 321560 305328 321612 305380
rect 321928 305328 321980 305380
rect 323216 305328 323268 305380
rect 323768 305328 323820 305380
rect 324412 305328 324464 305380
rect 325148 305328 325200 305380
rect 325976 305328 326028 305380
rect 326344 305328 326396 305380
rect 328644 305328 328696 305380
rect 329012 305328 329064 305380
rect 330208 305328 330260 305380
rect 331128 305328 331180 305380
rect 305092 305260 305144 305312
rect 305920 305260 305972 305312
rect 308128 305260 308180 305312
rect 308956 305260 309008 305312
rect 309232 305260 309284 305312
rect 309508 305260 309560 305312
rect 314752 305260 314804 305312
rect 315488 305260 315540 305312
rect 323032 305260 323084 305312
rect 323952 305260 324004 305312
rect 326068 305260 326120 305312
rect 326988 305260 327040 305312
rect 328736 305260 328788 305312
rect 329380 305260 329432 305312
rect 330116 305260 330168 305312
rect 330944 305260 330996 305312
rect 306380 305192 306432 305244
rect 307300 305192 307352 305244
rect 310520 305192 310572 305244
rect 311348 305192 311400 305244
rect 314660 305192 314712 305244
rect 315948 305192 316000 305244
rect 321560 305192 321612 305244
rect 322664 305192 322716 305244
rect 328552 305192 328604 305244
rect 329472 305192 329524 305244
rect 329932 305192 329984 305244
rect 330576 305192 330628 305244
rect 332508 305396 332560 305448
rect 338764 305396 338816 305448
rect 331404 305328 331456 305380
rect 332232 305328 332284 305380
rect 332784 305328 332836 305380
rect 333520 305328 333572 305380
rect 331956 305260 332008 305312
rect 339868 305260 339920 305312
rect 343640 305396 343692 305448
rect 254032 304784 254084 304836
rect 254308 304784 254360 304836
rect 254032 304648 254084 304700
rect 254492 304648 254544 304700
rect 316592 304444 316644 304496
rect 443644 304444 443696 304496
rect 85580 304376 85632 304428
rect 245660 304376 245712 304428
rect 319628 304376 319680 304428
rect 485044 304376 485096 304428
rect 82176 304308 82228 304360
rect 244372 304308 244424 304360
rect 325516 304308 325568 304360
rect 516784 304308 516836 304360
rect 7564 304240 7616 304292
rect 230480 304240 230532 304292
rect 233424 304240 233476 304292
rect 233608 304240 233660 304292
rect 256976 304240 257028 304292
rect 257252 304240 257304 304292
rect 276296 304240 276348 304292
rect 276572 304240 276624 304292
rect 304908 304240 304960 304292
rect 305460 304240 305512 304292
rect 310796 304240 310848 304292
rect 311164 304240 311216 304292
rect 313648 304240 313700 304292
rect 313924 304240 313976 304292
rect 318984 304240 319036 304292
rect 319260 304240 319312 304292
rect 334532 304240 334584 304292
rect 563704 304240 563756 304292
rect 291384 304172 291436 304224
rect 292304 304172 292356 304224
rect 230664 304104 230716 304156
rect 231768 304104 231820 304156
rect 248604 304104 248656 304156
rect 249616 304104 249668 304156
rect 251548 303968 251600 304020
rect 252468 303968 252520 304020
rect 273444 303968 273496 304020
rect 274272 303968 274324 304020
rect 318800 303696 318852 303748
rect 319904 303696 319956 303748
rect 275928 303560 275980 303612
rect 341248 303560 341300 303612
rect 272524 303492 272576 303544
rect 342352 303492 342404 303544
rect 264980 303424 265032 303476
rect 265900 303424 265952 303476
rect 272800 303424 272852 303476
rect 343732 303424 343784 303476
rect 269856 303356 269908 303408
rect 344836 303356 344888 303408
rect 279884 303288 279936 303340
rect 355140 303288 355192 303340
rect 269948 303220 270000 303272
rect 345112 303220 345164 303272
rect 270040 303152 270092 303204
rect 346400 303152 346452 303204
rect 278136 303084 278188 303136
rect 357532 303084 357584 303136
rect 93124 303016 93176 303068
rect 245108 303016 245160 303068
rect 276112 303016 276164 303068
rect 277216 303016 277268 303068
rect 278228 303016 278280 303068
rect 358912 303016 358964 303068
rect 93860 302948 93912 303000
rect 247224 302948 247276 303000
rect 275376 302948 275428 303000
rect 358820 302948 358872 303000
rect 8944 302880 8996 302932
rect 231400 302880 231452 302932
rect 275468 302880 275520 302932
rect 359096 302880 359148 302932
rect 277124 302812 277176 302864
rect 277308 302812 277360 302864
rect 293776 302812 293828 302864
rect 342812 302812 342864 302864
rect 263600 302744 263652 302796
rect 264612 302744 264664 302796
rect 294972 302744 295024 302796
rect 342536 302744 342588 302796
rect 293592 302676 293644 302728
rect 338120 302676 338172 302728
rect 258264 302608 258316 302660
rect 258540 302608 258592 302660
rect 320548 301588 320600 301640
rect 491944 301588 491996 301640
rect 48964 301520 49016 301572
rect 239128 301520 239180 301572
rect 328920 301520 328972 301572
rect 534724 301520 534776 301572
rect 43444 301452 43496 301504
rect 237380 301452 237432 301504
rect 334808 301452 334860 301504
rect 565820 301452 565872 301504
rect 285220 300772 285272 300824
rect 336924 300772 336976 300824
rect 285404 300704 285456 300756
rect 338304 300704 338356 300756
rect 290832 300636 290884 300688
rect 345020 300636 345072 300688
rect 286968 300568 287020 300620
rect 346584 300568 346636 300620
rect 267924 300500 267976 300552
rect 268292 300500 268344 300552
rect 296628 300500 296680 300552
rect 357624 300500 357676 300552
rect 241888 300432 241940 300484
rect 242072 300432 242124 300484
rect 283840 300432 283892 300484
rect 345296 300432 345348 300484
rect 282552 300364 282604 300416
rect 347320 300364 347372 300416
rect 285496 300296 285548 300348
rect 351092 300296 351144 300348
rect 292304 300228 292356 300280
rect 357900 300228 357952 300280
rect 53104 300160 53156 300212
rect 238852 300160 238904 300212
rect 279608 300160 279660 300212
rect 349344 300160 349396 300212
rect 10324 300092 10376 300144
rect 231032 300092 231084 300144
rect 285312 300092 285364 300144
rect 360200 300092 360252 300144
rect 286876 300024 286928 300076
rect 338212 300024 338264 300076
rect 288256 299956 288308 300008
rect 340512 299956 340564 300008
rect 290740 299888 290792 299940
rect 341432 299888 341484 299940
rect 313740 298936 313792 298988
rect 454040 298936 454092 298988
rect 323400 298868 323452 298920
rect 502984 298868 503036 298920
rect 326252 298800 326304 298852
rect 520280 298800 520332 298852
rect 53840 298732 53892 298784
rect 238760 298732 238812 298784
rect 333060 298732 333112 298784
rect 557540 298732 557592 298784
rect 251180 298596 251232 298648
rect 251364 298596 251416 298648
rect 278596 297780 278648 297832
rect 338396 297780 338448 297832
rect 282460 297712 282512 297764
rect 343824 297712 343876 297764
rect 275836 297644 275888 297696
rect 339684 297644 339736 297696
rect 283932 297576 283984 297628
rect 359004 297576 359056 297628
rect 323308 297508 323360 297560
rect 507860 297508 507912 297560
rect 86960 297440 87012 297492
rect 245936 297440 245988 297492
rect 269580 297440 269632 297492
rect 285864 297440 285916 297492
rect 332968 297440 333020 297492
rect 560300 297440 560352 297492
rect 60740 297372 60792 297424
rect 240416 297372 240468 297424
rect 269580 297236 269632 297288
rect 334256 297372 334308 297424
rect 570604 297372 570656 297424
rect 285956 297236 286008 297288
rect 93952 296012 94004 296064
rect 247592 296012 247644 296064
rect 316316 296012 316368 296064
rect 467104 296012 467156 296064
rect 66904 295944 66956 295996
rect 241980 295944 242032 295996
rect 324688 295944 324740 295996
rect 514024 295944 514076 295996
rect 316224 294720 316276 294772
rect 471244 294720 471296 294772
rect 69020 294652 69072 294704
rect 241796 294652 241848 294704
rect 327540 294652 327592 294704
rect 529940 294652 529992 294704
rect 31024 294584 31076 294636
rect 234896 294584 234948 294636
rect 283104 294584 283156 294636
rect 283288 294584 283340 294636
rect 328828 294584 328880 294636
rect 535460 294584 535512 294636
rect 3332 293904 3384 293956
rect 228456 293904 228508 293956
rect 54484 293224 54536 293276
rect 239036 293224 239088 293276
rect 327448 293224 327500 293276
rect 527824 293224 527876 293276
rect 71780 291864 71832 291916
rect 243084 291864 243136 291916
rect 34520 291796 34572 291848
rect 236276 291796 236328 291848
rect 328736 291796 328788 291848
rect 538864 291796 538916 291848
rect 269488 291116 269540 291168
rect 269672 291116 269724 291168
rect 331680 290504 331732 290556
rect 549904 290504 549956 290556
rect 41420 290436 41472 290488
rect 237656 290436 237708 290488
rect 334164 290436 334216 290488
rect 567200 290436 567252 290488
rect 58624 289144 58676 289196
rect 240324 289144 240376 289196
rect 331588 289144 331640 289196
rect 552664 289144 552716 289196
rect 13084 289076 13136 289128
rect 232136 289076 232188 289128
rect 334072 289076 334124 289128
rect 567844 289076 567896 289128
rect 312176 287784 312228 287836
rect 448520 287784 448572 287836
rect 312268 287716 312320 287768
rect 449900 287716 449952 287768
rect 9680 287648 9732 287700
rect 230664 287648 230716 287700
rect 332876 287648 332928 287700
rect 561680 287648 561732 287700
rect 315120 286492 315172 286544
rect 462320 286492 462372 286544
rect 318156 286424 318208 286476
rect 467840 286424 467892 286476
rect 89720 286356 89772 286408
rect 245844 286356 245896 286408
rect 319168 286356 319220 286408
rect 481640 286356 481692 286408
rect 46296 286288 46348 286340
rect 237564 286288 237616 286340
rect 335820 286288 335872 286340
rect 575480 286288 575532 286340
rect 96620 284996 96672 285048
rect 247316 284996 247368 285048
rect 39396 284928 39448 284980
rect 236184 284928 236236 284980
rect 313648 284928 313700 284980
rect 453304 284928 453356 284980
rect 313556 283704 313608 283756
rect 456800 283704 456852 283756
rect 67640 283636 67692 283688
rect 241704 283636 241756 283688
rect 317696 283636 317748 283688
rect 481732 283636 481784 283688
rect 16580 283568 16632 283620
rect 232044 283568 232096 283620
rect 333980 283568 334032 283620
rect 571340 283568 571392 283620
rect 318064 282276 318116 282328
rect 460940 282276 460992 282328
rect 74540 282208 74592 282260
rect 235264 282208 235316 282260
rect 315028 282208 315080 282260
rect 459560 282208 459612 282260
rect 20720 282140 20772 282192
rect 233608 282140 233660 282192
rect 319076 282140 319128 282192
rect 484400 282140 484452 282192
rect 320824 280916 320876 280968
rect 474740 280916 474792 280968
rect 88984 280848 89036 280900
rect 245752 280848 245804 280900
rect 316132 280848 316184 280900
rect 472624 280848 472676 280900
rect 26240 280780 26292 280832
rect 234804 280780 234856 280832
rect 321836 280780 321888 280832
rect 502340 280780 502392 280832
rect 92480 279488 92532 279540
rect 247224 279488 247276 279540
rect 318984 279488 319036 279540
rect 485780 279488 485832 279540
rect 40684 279420 40736 279472
rect 234712 279420 234764 279472
rect 324596 279420 324648 279472
rect 511264 279420 511316 279472
rect 317604 278128 317656 278180
rect 477500 278128 477552 278180
rect 323216 278060 323268 278112
rect 509240 278060 509292 278112
rect 35164 277992 35216 278044
rect 236092 277992 236144 278044
rect 330392 277992 330444 278044
rect 542360 277992 542412 278044
rect 310796 276700 310848 276752
rect 440240 276700 440292 276752
rect 35900 276632 35952 276684
rect 236368 276632 236420 276684
rect 320456 276632 320508 276684
rect 496084 276632 496136 276684
rect 310704 275408 310756 275460
rect 444380 275408 444432 275460
rect 44180 275340 44232 275392
rect 236736 275340 236788 275392
rect 321744 275340 321796 275392
rect 499580 275340 499632 275392
rect 22744 275272 22796 275324
rect 233516 275272 233568 275324
rect 327356 275272 327408 275324
rect 531320 275272 531372 275324
rect 312084 274116 312136 274168
rect 448612 274116 448664 274168
rect 323124 274048 323176 274100
rect 506480 274048 506532 274100
rect 14464 273980 14516 274032
rect 230940 273980 230992 274032
rect 328644 273980 328696 274032
rect 536104 273980 536156 274032
rect 99288 273912 99340 273964
rect 336832 273912 336884 273964
rect 367744 273164 367796 273216
rect 579896 273164 579948 273216
rect 326160 272552 326212 272604
rect 521660 272552 521712 272604
rect 50344 272484 50396 272536
rect 238944 272484 238996 272536
rect 332784 272484 332836 272536
rect 560944 272484 560996 272536
rect 311992 271192 312044 271244
rect 450544 271192 450596 271244
rect 52460 271124 52512 271176
rect 239312 271124 239364 271176
rect 328552 271124 328604 271176
rect 540244 271124 540296 271176
rect 313464 269900 313516 269952
rect 458180 269900 458232 269952
rect 327264 269832 327316 269884
rect 528560 269832 528612 269884
rect 57336 269764 57388 269816
rect 240232 269764 240284 269816
rect 331496 269764 331548 269816
rect 552020 269764 552072 269816
rect 314936 268472 314988 268524
rect 464344 268472 464396 268524
rect 328460 268404 328512 268456
rect 539692 268404 539744 268456
rect 59360 268336 59412 268388
rect 240508 268336 240560 268388
rect 331404 268336 331456 268388
rect 556252 268336 556304 268388
rect 2964 267656 3016 267708
rect 224224 267656 224276 267708
rect 238300 267112 238352 267164
rect 350816 267112 350868 267164
rect 317512 267044 317564 267096
rect 476120 267044 476172 267096
rect 332692 266976 332744 267028
rect 558920 266976 558972 267028
rect 318892 265752 318944 265804
rect 488540 265752 488592 265804
rect 331312 265684 331364 265736
rect 554044 265684 554096 265736
rect 62120 265616 62172 265668
rect 241612 265616 241664 265668
rect 335728 265616 335780 265668
rect 574744 265616 574796 265668
rect 309600 264392 309652 264444
rect 436744 264392 436796 264444
rect 310612 264324 310664 264376
rect 440332 264324 440384 264376
rect 314844 264256 314896 264308
rect 463700 264256 463752 264308
rect 66260 264188 66312 264240
rect 241888 264188 241940 264240
rect 320364 264188 320416 264240
rect 491300 264188 491352 264240
rect 238392 263032 238444 263084
rect 360384 263032 360436 263084
rect 314752 262964 314804 263016
rect 456064 262964 456116 263016
rect 75184 262896 75236 262948
rect 243268 262896 243320 262948
rect 318800 262896 318852 262948
rect 490012 262896 490064 262948
rect 4160 262828 4212 262880
rect 229744 262828 229796 262880
rect 320272 262828 320324 262880
rect 495440 262828 495492 262880
rect 320180 261604 320232 261656
rect 492680 261604 492732 261656
rect 77300 261536 77352 261588
rect 243176 261536 243228 261588
rect 321652 261536 321704 261588
rect 494796 261536 494848 261588
rect 21364 261468 21416 261520
rect 233424 261468 233476 261520
rect 330300 261468 330352 261520
rect 546500 261468 546552 261520
rect 364984 260176 365036 260228
rect 580448 260176 580500 260228
rect 42800 260108 42852 260160
rect 237472 260108 237524 260160
rect 330208 260108 330260 260160
rect 549260 260108 549312 260160
rect 91100 258748 91152 258800
rect 246028 258748 246080 258800
rect 313372 258748 313424 258800
rect 452660 258748 452712 258800
rect 13820 258680 13872 258732
rect 231952 258680 232004 258732
rect 363604 258680 363656 258732
rect 580356 258680 580408 258732
rect 326068 257388 326120 257440
rect 527180 257388 527232 257440
rect 373264 257320 373316 257372
rect 581092 257320 581144 257372
rect 325976 255960 326028 256012
rect 523040 255960 523092 256012
rect 3148 255212 3200 255264
rect 220084 255212 220136 255264
rect 316040 254668 316092 254720
rect 471980 254668 472032 254720
rect 317420 254600 317472 254652
rect 478144 254600 478196 254652
rect 88340 254532 88392 254584
rect 236644 254532 236696 254584
rect 330116 254532 330168 254584
rect 547880 254532 547932 254584
rect 297732 253308 297784 253360
rect 335636 253308 335688 253360
rect 98000 253240 98052 253292
rect 247500 253240 247552 253292
rect 335452 253240 335504 253292
rect 574100 253240 574152 253292
rect 30380 253172 30432 253224
rect 234988 253172 235040 253224
rect 335544 253172 335596 253224
rect 578240 253172 578292 253224
rect 297272 252016 297324 252068
rect 344008 252016 344060 252068
rect 323032 251948 323084 252000
rect 510620 251948 510672 252000
rect 324504 251880 324556 251932
rect 514116 251880 514168 251932
rect 17960 251812 18012 251864
rect 233332 251812 233384 251864
rect 332600 251812 332652 251864
rect 564532 251812 564584 251864
rect 238484 250724 238536 250776
rect 356336 250724 356388 250776
rect 359372 250724 359424 250776
rect 441712 250724 441764 250776
rect 310520 250656 310572 250708
rect 441620 250656 441672 250708
rect 311900 250588 311952 250640
rect 445760 250588 445812 250640
rect 321560 250520 321612 250572
rect 503720 250520 503772 250572
rect 22100 250452 22152 250504
rect 233700 250452 233752 250504
rect 330024 250452 330076 250504
rect 545120 250452 545172 250504
rect 313280 249160 313332 249212
rect 456892 249160 456944 249212
rect 314660 249092 314712 249144
rect 466460 249092 466512 249144
rect 12440 249024 12492 249076
rect 232228 249024 232280 249076
rect 335360 249024 335412 249076
rect 571984 249024 572036 249076
rect 298836 248344 298888 248396
rect 347964 248344 348016 248396
rect 360292 248344 360344 248396
rect 438216 248344 438268 248396
rect 292488 248276 292540 248328
rect 345204 248276 345256 248328
rect 356244 248276 356296 248328
rect 436928 248276 436980 248328
rect 297824 248208 297876 248260
rect 350724 248208 350776 248260
rect 359280 248208 359332 248260
rect 441804 248208 441856 248260
rect 286692 248140 286744 248192
rect 346676 248140 346728 248192
rect 357808 248140 357860 248192
rect 440608 248140 440660 248192
rect 288164 248072 288216 248124
rect 348240 248072 348292 248124
rect 357716 248072 357768 248124
rect 441896 248072 441948 248124
rect 288072 248004 288124 248056
rect 305460 248004 305512 248056
rect 306932 248004 306984 248056
rect 437480 248004 437532 248056
rect 289176 247936 289228 247988
rect 303896 247936 303948 247988
rect 308220 247936 308272 247988
rect 438860 247936 438912 247988
rect 290648 247868 290700 247920
rect 305184 247868 305236 247920
rect 309508 247868 309560 247920
rect 440424 247868 440476 247920
rect 292396 247800 292448 247852
rect 305368 247800 305420 247852
rect 322940 247800 322992 247852
rect 506572 247800 506624 247852
rect 324412 247732 324464 247784
rect 517520 247732 517572 247784
rect 4804 247664 4856 247716
rect 229192 247664 229244 247716
rect 287888 247664 287940 247716
rect 300676 247664 300728 247716
rect 329932 247664 329984 247716
rect 547972 247664 548024 247716
rect 300768 247596 300820 247648
rect 346768 247596 346820 247648
rect 297088 247528 297140 247580
rect 339592 247528 339644 247580
rect 288992 247460 289044 247512
rect 303804 247460 303856 247512
rect 286784 247392 286836 247444
rect 303988 247392 304040 247444
rect 298744 247052 298796 247104
rect 304080 247052 304132 247104
rect 297364 246984 297416 247036
rect 342720 246984 342772 247036
rect 298928 246916 298980 246968
rect 345480 246916 345532 246968
rect 299388 246848 299440 246900
rect 351000 246848 351052 246900
rect 297180 246780 297232 246832
rect 349436 246780 349488 246832
rect 296536 246712 296588 246764
rect 350908 246712 350960 246764
rect 289636 246644 289688 246696
rect 349252 246644 349304 246696
rect 325884 246576 325936 246628
rect 524420 246576 524472 246628
rect 325792 246508 325844 246560
rect 525800 246508 525852 246560
rect 327172 246440 327224 246492
rect 534080 246440 534132 246492
rect 329840 246372 329892 246424
rect 543740 246372 543792 246424
rect 3608 246304 3660 246356
rect 228364 246304 228416 246356
rect 331220 246304 331272 246356
rect 553400 246304 553452 246356
rect 297456 246236 297508 246288
rect 341156 246236 341208 246288
rect 291016 245556 291068 245608
rect 306656 245556 306708 245608
rect 309416 245556 309468 245608
rect 437940 245556 437992 245608
rect 292212 245488 292264 245540
rect 305092 245488 305144 245540
rect 307944 245488 307996 245540
rect 437664 245488 437716 245540
rect 293684 245420 293736 245472
rect 303712 245420 303764 245472
rect 309324 245420 309376 245472
rect 439136 245420 439188 245472
rect 293408 245352 293460 245404
rect 303620 245352 303672 245404
rect 307852 245352 307904 245404
rect 437848 245352 437900 245404
rect 295248 245284 295300 245336
rect 305000 245284 305052 245336
rect 309140 245284 309192 245336
rect 439320 245284 439372 245336
rect 306840 245216 306892 245268
rect 437572 245216 437624 245268
rect 295156 245148 295208 245200
rect 300860 245148 300912 245200
rect 306472 245148 306524 245200
rect 437756 245148 437808 245200
rect 292488 245080 292540 245132
rect 299572 245080 299624 245132
rect 308036 245080 308088 245132
rect 439412 245080 439464 245132
rect 291108 245012 291160 245064
rect 299664 245012 299716 245064
rect 307760 245012 307812 245064
rect 439228 245012 439280 245064
rect 291016 244944 291068 244996
rect 301136 244944 301188 244996
rect 306748 244944 306800 244996
rect 438952 244944 439004 244996
rect 7656 244876 7708 244928
rect 230848 244876 230900 244928
rect 289728 244876 289780 244928
rect 302240 244876 302292 244928
rect 306380 244876 306432 244928
rect 439044 244876 439096 244928
rect 299112 244808 299164 244860
rect 342628 244808 342680 244860
rect 356520 244808 356572 244860
rect 438308 244808 438360 244860
rect 299020 244740 299072 244792
rect 339776 244740 339828 244792
rect 360476 244740 360528 244792
rect 439688 244740 439740 244792
rect 297640 244672 297692 244724
rect 337016 244672 337068 244724
rect 295248 244604 295300 244656
rect 299480 244604 299532 244656
rect 288348 244468 288400 244520
rect 291752 244468 291804 244520
rect 291752 244332 291804 244384
rect 299296 244332 299348 244384
rect 293684 243720 293736 243772
rect 300768 243720 300820 243772
rect 299296 243652 299348 243704
rect 343916 243652 343968 243704
rect 299204 243584 299256 243636
rect 345388 243584 345440 243636
rect 97816 243516 97868 243568
rect 297272 243516 297324 243568
rect 297916 243516 297968 243568
rect 356060 243516 356112 243568
rect 97908 243448 97960 243500
rect 298744 243448 298796 243500
rect 299020 243448 299072 243500
rect 97724 243380 97776 243432
rect 298928 243380 298980 243432
rect 3240 241408 3292 241460
rect 98644 241408 98696 241460
rect 3332 215228 3384 215280
rect 86224 215228 86276 215280
rect 292212 198024 292264 198076
rect 297180 198024 297232 198076
rect 297548 197412 297600 197464
rect 298836 197412 298888 197464
rect 292396 197276 292448 197328
rect 298836 197276 298888 197328
rect 296628 195916 296680 195968
rect 298376 195916 298428 195968
rect 3148 188980 3200 189032
rect 95976 188980 96028 189032
rect 261116 177284 261168 177336
rect 277676 177284 277728 177336
rect 285220 171028 285272 171080
rect 297180 171028 297232 171080
rect 236736 170348 236788 170400
rect 285220 170348 285272 170400
rect 238576 167628 238628 167680
rect 297732 167628 297784 167680
rect 292304 166948 292356 167000
rect 296720 166948 296772 167000
rect 3516 164160 3568 164212
rect 84844 164160 84896 164212
rect 97816 159876 97868 159928
rect 298928 159876 298980 159928
rect 97632 159808 97684 159860
rect 297272 159808 297324 159860
rect 97540 159740 97592 159792
rect 297364 159740 297416 159792
rect 97448 159672 97500 159724
rect 238576 159672 238628 159724
rect 97908 159604 97960 159656
rect 236736 159604 236788 159656
rect 284484 159604 284536 159656
rect 299480 159604 299532 159656
rect 287612 159536 287664 159588
rect 309140 159536 309192 159588
rect 293316 159468 293368 159520
rect 327172 159468 327224 159520
rect 234620 159400 234672 159452
rect 273720 159400 273772 159452
rect 298192 159400 298244 159452
rect 338764 159400 338816 159452
rect 220820 159332 220872 159384
rect 271052 159332 271104 159384
rect 298836 159332 298888 159384
rect 348240 159332 348292 159384
rect 293684 159264 293736 159316
rect 351000 159264 351052 159316
rect 297548 159196 297600 159248
rect 356060 159196 356112 159248
rect 286784 159128 286836 159180
rect 353576 159128 353628 159180
rect 165988 159060 166040 159112
rect 238116 159060 238168 159112
rect 299388 159060 299440 159112
rect 368296 159060 368348 159112
rect 160928 158992 160980 159044
rect 240784 158992 240836 159044
rect 296536 158992 296588 159044
rect 365904 158992 365956 159044
rect 156052 158924 156104 158976
rect 249064 158924 249116 158976
rect 288164 158924 288216 158976
rect 358452 158924 358504 158976
rect 153660 158856 153712 158908
rect 250536 158856 250588 158908
rect 289636 158856 289688 158908
rect 360936 158856 360988 158908
rect 168288 158788 168340 158840
rect 286416 158788 286468 158840
rect 292212 158788 292264 158840
rect 363420 158788 363472 158840
rect 175924 158720 175976 158772
rect 296168 158720 296220 158772
rect 297824 158720 297876 158772
rect 370964 158720 371016 158772
rect 388536 158720 388588 158772
rect 436928 158720 436980 158772
rect 128728 158652 128780 158704
rect 276020 158652 276072 158704
rect 293776 158652 293828 158704
rect 338396 158652 338448 158704
rect 373448 158652 373500 158704
rect 440516 158652 440568 158704
rect 126520 158584 126572 158636
rect 276572 158584 276624 158636
rect 276848 158584 276900 158636
rect 298008 158584 298060 158636
rect 331220 158584 331272 158636
rect 376024 158584 376076 158636
rect 438124 158584 438176 158636
rect 121920 158516 121972 158568
rect 290740 158516 290792 158568
rect 294972 158516 295024 158568
rect 340972 158516 341024 158568
rect 378600 158516 378652 158568
rect 439596 158516 439648 158568
rect 120632 158448 120684 158500
rect 288256 158448 288308 158500
rect 290648 158448 290700 158500
rect 290924 158448 290976 158500
rect 293592 158448 293644 158500
rect 328276 158448 328328 158500
rect 380992 158448 381044 158500
rect 436836 158448 436888 158500
rect 282460 158380 282512 158432
rect 343548 158380 343600 158432
rect 383568 158380 383620 158432
rect 438032 158380 438084 158432
rect 127624 158312 127676 158364
rect 295064 158312 295116 158364
rect 327540 158312 327592 158364
rect 385960 158312 386012 158364
rect 439504 158312 439556 158364
rect 132408 158244 132460 158296
rect 299204 158244 299256 158296
rect 332324 158244 332376 158296
rect 391480 158244 391532 158296
rect 438308 158244 438360 158296
rect 131304 158176 131356 158228
rect 298008 158176 298060 158228
rect 299388 158176 299440 158228
rect 329932 158176 329984 158228
rect 394240 158176 394292 158228
rect 440608 158176 440660 158228
rect 275928 158108 275980 158160
rect 336004 158108 336056 158160
rect 395896 158108 395948 158160
rect 441896 158108 441948 158160
rect 133512 158040 133564 158092
rect 283840 158040 283892 158092
rect 286140 158040 286192 158092
rect 286876 158040 286928 158092
rect 319444 158040 319496 158092
rect 398472 158040 398524 158092
rect 441712 158040 441764 158092
rect 275836 157972 275888 158024
rect 333612 157972 333664 158024
rect 401048 157972 401100 158024
rect 441804 157972 441856 158024
rect 159640 157904 159692 157956
rect 285128 157904 285180 157956
rect 288256 157904 288308 157956
rect 320548 157904 320600 157956
rect 403992 157904 404044 157956
rect 438216 157904 438268 157956
rect 188712 157836 188764 157888
rect 238484 157836 238536 157888
rect 290740 157836 290792 157888
rect 321652 157836 321704 157888
rect 406476 157836 406528 157888
rect 439688 157836 439740 157888
rect 206008 157768 206060 157820
rect 238392 157768 238444 157820
rect 119896 157700 119948 157752
rect 286140 157700 286192 157752
rect 97724 157632 97776 157684
rect 297456 157632 297508 157684
rect 130568 157564 130620 157616
rect 299388 157564 299440 157616
rect 331312 157496 331364 157548
rect 354404 157496 354456 157548
rect 329748 157428 329800 157480
rect 356980 157428 357032 157480
rect 327264 157360 327316 157412
rect 355232 157360 355284 157412
rect 116216 157292 116268 157344
rect 283748 157292 283800 157344
rect 284024 157292 284076 157344
rect 284484 157292 284536 157344
rect 285588 157292 285640 157344
rect 347596 157292 347648 157344
rect 118240 157224 118292 157276
rect 285404 157224 285456 157276
rect 290924 157224 290976 157276
rect 135904 156952 135956 157004
rect 282552 157156 282604 157208
rect 335820 157156 335872 157208
rect 280068 157088 280120 157140
rect 339316 157088 339368 157140
rect 278596 157020 278648 157072
rect 330300 157020 330352 157072
rect 137008 156884 137060 156936
rect 282828 156952 282880 157004
rect 336924 156952 336976 157004
rect 286140 156884 286192 156936
rect 286968 156884 287020 156936
rect 334532 156884 334584 156936
rect 138388 156816 138440 156868
rect 279976 156816 280028 156868
rect 283748 156816 283800 156868
rect 316040 156816 316092 156868
rect 139676 156748 139728 156800
rect 280068 156748 280120 156800
rect 290648 156748 290700 156800
rect 323124 156748 323176 156800
rect 282920 156680 282972 156732
rect 284116 156680 284168 156732
rect 317052 156680 317104 156732
rect 125600 156612 125652 156664
rect 252836 156612 252888 156664
rect 253296 156612 253348 156664
rect 275008 156612 275060 156664
rect 290188 156612 290240 156664
rect 331220 156612 331272 156664
rect 184020 156544 184072 156596
rect 280988 156544 281040 156596
rect 287520 156544 287572 156596
rect 313280 156544 313332 156596
rect 185952 156476 186004 156528
rect 280896 156476 280948 156528
rect 285956 156476 286008 156528
rect 302240 156476 302292 156528
rect 191472 156408 191524 156460
rect 280804 156408 280856 156460
rect 279976 156340 280028 156392
rect 338120 156340 338172 156392
rect 123944 156272 123996 156324
rect 290648 156272 290700 156324
rect 134616 156204 134668 156256
rect 286140 156204 286192 156256
rect 117320 156136 117372 156188
rect 282920 156136 282972 156188
rect 148692 156068 148744 156120
rect 284484 156068 284536 156120
rect 271144 155864 271196 155916
rect 276388 155864 276440 155916
rect 283564 155864 283616 155916
rect 285956 155864 286008 155916
rect 286140 155864 286192 155916
rect 345112 155864 345164 155916
rect 276020 155796 276072 155848
rect 277216 155796 277268 155848
rect 346400 155796 346452 155848
rect 141792 155728 141844 155780
rect 285496 155728 285548 155780
rect 341156 155728 341208 155780
rect 282368 155660 282420 155712
rect 282644 155660 282696 155712
rect 348700 155660 348752 155712
rect 143080 155592 143132 155644
rect 282736 155592 282788 155644
rect 342352 155592 342404 155644
rect 140688 155524 140740 155576
rect 279608 155524 279660 155576
rect 339592 155524 339644 155576
rect 148784 155456 148836 155508
rect 282368 155456 282420 155508
rect 282920 155456 282972 155508
rect 284208 155456 284260 155508
rect 343916 155456 343968 155508
rect 145288 155388 145340 155440
rect 279700 155388 279752 155440
rect 286140 155388 286192 155440
rect 289544 155388 289596 155440
rect 324228 155388 324280 155440
rect 146392 155320 146444 155372
rect 276020 155320 276072 155372
rect 299388 155320 299440 155372
rect 327264 155320 327316 155372
rect 148416 155252 148468 155304
rect 269948 155252 270000 155304
rect 288900 155252 288952 155304
rect 320180 155252 320232 155304
rect 150992 155184 151044 155236
rect 270040 155184 270092 155236
rect 291660 155184 291712 155236
rect 338120 155184 338172 155236
rect 201040 155116 201092 155168
rect 275376 155116 275428 155168
rect 286048 155116 286100 155168
rect 306380 155116 306432 155168
rect 203432 155048 203484 155100
rect 275468 155048 275520 155100
rect 229100 154980 229152 155032
rect 272248 154980 272300 155032
rect 155776 154912 155828 154964
rect 298376 154912 298428 154964
rect 299388 154912 299440 154964
rect 124772 154844 124824 154896
rect 289544 154844 289596 154896
rect 144000 154776 144052 154828
rect 282920 154776 282972 154828
rect 125416 154504 125468 154556
rect 276020 154504 276072 154556
rect 279792 154504 279844 154556
rect 280068 154504 280120 154556
rect 351092 154504 351144 154556
rect 153844 154436 153896 154488
rect 297916 154436 297968 154488
rect 353300 154436 353352 154488
rect 152648 154368 152700 154420
rect 141516 154300 141568 154352
rect 272524 154300 272576 154352
rect 290832 154368 290884 154420
rect 345756 154368 345808 154420
rect 281356 154300 281408 154352
rect 352196 154300 352248 154352
rect 149888 154232 149940 154284
rect 279884 154232 279936 154284
rect 349804 154232 349856 154284
rect 276020 154164 276072 154216
rect 277308 154164 277360 154216
rect 324872 154164 324924 154216
rect 151360 154096 151412 154148
rect 280068 154096 280120 154148
rect 157064 154028 157116 154080
rect 283932 154028 283984 154080
rect 329748 154096 329800 154148
rect 297456 154028 297508 154080
rect 331312 154028 331364 154080
rect 146024 153960 146076 154012
rect 269856 153960 269908 154012
rect 195888 153892 195940 153944
rect 278136 153892 278188 153944
rect 164240 153824 164292 153876
rect 259920 153824 259972 153876
rect 287428 153824 287480 153876
rect 316040 153824 316092 153876
rect 198464 153756 198516 153808
rect 278228 153756 278280 153808
rect 202880 153688 202932 153740
rect 266820 153688 266872 153740
rect 231860 153620 231912 153672
rect 272156 153620 272208 153672
rect 154488 153552 154540 153604
rect 296720 153552 296772 153604
rect 297456 153552 297508 153604
rect 233240 152668 233292 152720
rect 272064 152668 272116 152720
rect 227720 152600 227772 152652
rect 269764 152600 269816 152652
rect 288808 152600 288860 152652
rect 324320 152600 324372 152652
rect 193220 152532 193272 152584
rect 265440 152532 265492 152584
rect 294328 152532 294380 152584
rect 349160 152532 349212 152584
rect 168380 152464 168432 152516
rect 242256 152464 242308 152516
rect 299112 152464 299164 152516
rect 376760 152464 376812 152516
rect 272524 151784 272576 151836
rect 278964 151784 279016 151836
rect 209780 151172 209832 151224
rect 268108 151172 268160 151224
rect 284392 151172 284444 151224
rect 299572 151172 299624 151224
rect 175280 151104 175332 151156
rect 261484 151104 261536 151156
rect 290096 151104 290148 151156
rect 324412 151104 324464 151156
rect 146300 151036 146352 151088
rect 257160 151036 257212 151088
rect 292948 151036 293000 151088
rect 340880 151036 340932 151088
rect 268200 150424 268252 150476
rect 273904 150424 273956 150476
rect 213920 149812 213972 149864
rect 269580 149812 269632 149864
rect 285864 149812 285916 149864
rect 303620 149812 303672 149864
rect 184940 149744 184992 149796
rect 264060 149744 264112 149796
rect 292856 149744 292908 149796
rect 345020 149744 345072 149796
rect 157340 149676 157392 149728
rect 258356 149676 258408 149728
rect 295708 149676 295760 149728
rect 357440 149676 357492 149728
rect 215300 148452 215352 148504
rect 269488 148452 269540 148504
rect 189080 148384 189132 148436
rect 263968 148384 264020 148436
rect 291568 148384 291620 148436
rect 332600 148384 332652 148436
rect 135260 148316 135312 148368
rect 254216 148316 254268 148368
rect 294236 148316 294288 148368
rect 351920 148316 351972 148368
rect 176660 146956 176712 147008
rect 262496 146956 262548 147008
rect 287336 146956 287388 147008
rect 310520 146956 310572 147008
rect 128360 146888 128412 146940
rect 252744 146888 252796 146940
rect 253388 146888 253440 146940
rect 273628 146888 273680 146940
rect 290004 146888 290056 146940
rect 328460 146888 328512 146940
rect 279516 146548 279568 146600
rect 280436 146548 280488 146600
rect 219440 145664 219492 145716
rect 270868 145664 270920 145716
rect 287244 145664 287296 145716
rect 314660 145664 314712 145716
rect 195980 145596 196032 145648
rect 265348 145596 265400 145648
rect 292764 145596 292816 145648
rect 342260 145596 342312 145648
rect 153200 145528 153252 145580
rect 255964 145528 256016 145580
rect 265624 145528 265676 145580
rect 274916 145528 274968 145580
rect 275008 145528 275060 145580
rect 280344 145528 280396 145580
rect 283196 145528 283248 145580
rect 287244 145528 287296 145580
rect 294144 145528 294196 145580
rect 350540 145528 350592 145580
rect 218060 144304 218112 144356
rect 269396 144304 269448 144356
rect 154580 144236 154632 144288
rect 258264 144236 258316 144288
rect 288716 144236 288768 144288
rect 317420 144236 317472 144288
rect 143540 144168 143592 144220
rect 255780 144168 255832 144220
rect 294052 144168 294104 144220
rect 353300 144168 353352 144220
rect 269764 144032 269816 144084
rect 276296 144032 276348 144084
rect 236000 142944 236052 142996
rect 273536 142944 273588 142996
rect 183560 142876 183612 142928
rect 263876 142876 263928 142928
rect 288624 142876 288676 142928
rect 321560 142876 321612 142928
rect 132500 142808 132552 142860
rect 253204 142808 253256 142860
rect 295616 142808 295668 142860
rect 360200 142808 360252 142860
rect 193312 141516 193364 141568
rect 265256 141516 265308 141568
rect 139400 141448 139452 141500
rect 254584 141448 254636 141500
rect 285772 141448 285824 141500
rect 305000 141448 305052 141500
rect 121460 141380 121512 141432
rect 251548 141380 251600 141432
rect 291476 141380 291528 141432
rect 335360 141380 335412 141432
rect 197360 140156 197412 140208
rect 266728 140156 266780 140208
rect 285036 140156 285088 140208
rect 291476 140156 291528 140208
rect 150440 140088 150492 140140
rect 257068 140088 257120 140140
rect 114560 140020 114612 140072
rect 243636 140020 243688 140072
rect 291384 140020 291436 140072
rect 339500 140020 339552 140072
rect 201500 138728 201552 138780
rect 266636 138728 266688 138780
rect 126980 138660 127032 138712
rect 252652 138660 252704 138712
rect 292672 138660 292724 138712
rect 346400 138660 346452 138712
rect 3516 137912 3568 137964
rect 80704 137912 80756 137964
rect 211160 137368 211212 137420
rect 268016 137368 268068 137420
rect 161480 137300 161532 137352
rect 259828 137300 259880 137352
rect 107660 137232 107712 137284
rect 246488 137232 246540 137284
rect 293960 137232 294012 137284
rect 349252 137232 349304 137284
rect 222200 136008 222252 136060
rect 270776 136008 270828 136060
rect 165620 135940 165672 135992
rect 259736 135940 259788 135992
rect 103520 135872 103572 135924
rect 248696 135872 248748 135924
rect 168472 134580 168524 134632
rect 261300 134580 261352 134632
rect 147680 134512 147732 134564
rect 256976 134512 257028 134564
rect 288532 134512 288584 134564
rect 318800 134512 318852 134564
rect 191840 133220 191892 133272
rect 265164 133220 265216 133272
rect 172520 133152 172572 133204
rect 261208 133152 261260 133204
rect 261484 133152 261536 133204
rect 276204 133152 276256 133204
rect 216680 131860 216732 131912
rect 269304 131860 269356 131912
rect 179420 131792 179472 131844
rect 262404 131792 262456 131844
rect 110420 131724 110472 131776
rect 249984 131724 250036 131776
rect 288440 131724 288492 131776
rect 322940 131724 322992 131776
rect 230480 130500 230532 130552
rect 271972 130500 272024 130552
rect 186320 130432 186372 130484
rect 263784 130432 263836 130484
rect 100760 130364 100812 130416
rect 247776 130364 247828 130416
rect 289912 130364 289964 130416
rect 325700 130364 325752 130416
rect 190460 129072 190512 129124
rect 265072 129072 265124 129124
rect 149060 129004 149112 129056
rect 256884 129004 256936 129056
rect 291292 129004 291344 129056
rect 332692 129004 332744 129056
rect 204260 127644 204312 127696
rect 266544 127644 266596 127696
rect 131120 127576 131172 127628
rect 254124 127576 254176 127628
rect 291200 127576 291252 127628
rect 336740 127576 336792 127628
rect 208400 126284 208452 126336
rect 267924 126284 267976 126336
rect 138020 126216 138072 126268
rect 255688 126216 255740 126268
rect 294604 126216 294656 126268
rect 340972 126216 341024 126268
rect 280344 125536 280396 125588
rect 281908 125536 281960 125588
rect 218152 124924 218204 124976
rect 269212 124924 269264 124976
rect 169760 124856 169812 124908
rect 261024 124856 261076 124908
rect 269856 124856 269908 124908
rect 277584 124856 277636 124908
rect 296076 124856 296128 124908
rect 354680 124856 354732 124908
rect 278136 124448 278188 124500
rect 280252 124448 280304 124500
rect 226340 123496 226392 123548
rect 270684 123496 270736 123548
rect 158720 123428 158772 123480
rect 258172 123428 258224 123480
rect 133880 122068 133932 122120
rect 254032 122068 254084 122120
rect 254584 122068 254636 122120
rect 274824 122068 274876 122120
rect 136640 120708 136692 120760
rect 255596 120708 255648 120760
rect 140780 119348 140832 119400
rect 255504 119348 255556 119400
rect 151912 117920 151964 117972
rect 256792 117920 256844 117972
rect 143632 116560 143684 116612
rect 255412 116560 255464 116612
rect 127072 115200 127124 115252
rect 252928 115200 252980 115252
rect 162860 113772 162912 113824
rect 259644 113772 259696 113824
rect 460204 113092 460256 113144
rect 579804 113092 579856 113144
rect 167000 112412 167052 112464
rect 259552 112412 259604 112464
rect 3148 111732 3200 111784
rect 82084 111732 82136 111784
rect 173900 111052 173952 111104
rect 260932 111052 260984 111104
rect 180800 109692 180852 109744
rect 262312 109692 262364 109744
rect 185032 108264 185084 108316
rect 263692 108264 263744 108316
rect 198740 106904 198792 106956
rect 266452 106904 266504 106956
rect 187700 105544 187752 105596
rect 263600 105544 263652 105596
rect 205640 104116 205692 104168
rect 267832 104116 267884 104168
rect 223580 102824 223632 102876
rect 270592 102824 270644 102876
rect 118700 102756 118752 102808
rect 251456 102756 251508 102808
rect 135352 101396 135404 101448
rect 254400 101396 254452 101448
rect 234712 99968 234764 100020
rect 272340 99968 272392 100020
rect 144920 98608 144972 98660
rect 256700 98608 256752 98660
rect 3516 97928 3568 97980
rect 57244 97928 57296 97980
rect 155960 97248 156012 97300
rect 258540 97248 258592 97300
rect 111800 94460 111852 94512
rect 249892 94460 249944 94512
rect 115940 93100 115992 93152
rect 251364 93100 251416 93152
rect 106280 91740 106332 91792
rect 248604 91740 248656 91792
rect 99380 90312 99432 90364
rect 247408 90312 247460 90364
rect 49700 88952 49752 89004
rect 239220 88952 239272 89004
rect 117320 87592 117372 87644
rect 251272 87592 251324 87644
rect 113180 86232 113232 86284
rect 250076 86232 250128 86284
rect 3516 85484 3568 85536
rect 79324 85484 79376 85536
rect 446404 73108 446456 73160
rect 580172 73108 580224 73160
rect 142160 54476 142212 54528
rect 255872 54476 255924 54528
rect 194600 53048 194652 53100
rect 264980 53048 265032 53100
rect 494704 33056 494756 33108
rect 580172 33056 580224 33108
rect 47584 32376 47636 32428
rect 237748 32376 237800 32428
rect 295984 29588 296036 29640
rect 347780 29588 347832 29640
rect 110512 24080 110564 24132
rect 246396 24080 246448 24132
rect 102140 22720 102192 22772
rect 246304 22720 246356 22772
rect 212540 21360 212592 21412
rect 269120 21360 269172 21412
rect 209872 19932 209924 19984
rect 267740 19932 267792 19984
rect 201592 18572 201644 18624
rect 266912 18572 266964 18624
rect 160192 17280 160244 17332
rect 260012 17280 260064 17332
rect 259552 17212 259604 17264
rect 277492 17212 277544 17264
rect 292580 17212 292632 17264
rect 343640 17212 343692 17264
rect 177856 15852 177908 15904
rect 262680 15852 262732 15904
rect 289820 15852 289872 15904
rect 330392 15852 330444 15904
rect 120632 14424 120684 14476
rect 247684 14424 247736 14476
rect 264152 14424 264204 14476
rect 277400 14424 277452 14476
rect 287152 14424 287204 14476
rect 312176 14424 312228 14476
rect 260196 13132 260248 13184
rect 276112 13132 276164 13184
rect 123024 13064 123076 13116
rect 250444 13064 250496 13116
rect 276020 13064 276072 13116
rect 280528 13064 280580 13116
rect 285680 13064 285732 13116
rect 307944 13064 307996 13116
rect 255872 12452 255924 12504
rect 257344 12452 257396 12504
rect 160100 11772 160152 11824
rect 161296 11772 161348 11824
rect 184940 11772 184992 11824
rect 186136 11772 186188 11824
rect 234620 11772 234672 11824
rect 235816 11772 235868 11824
rect 284944 11772 284996 11824
rect 293224 11772 293276 11824
rect 105728 11704 105780 11756
rect 248512 11704 248564 11756
rect 266544 11704 266596 11756
rect 278044 11704 278096 11756
rect 287060 11704 287112 11756
rect 316224 11704 316276 11756
rect 272432 10480 272484 10532
rect 279332 10480 279384 10532
rect 60832 10276 60884 10328
rect 239404 10276 239456 10328
rect 244648 10276 244700 10328
rect 274732 10276 274784 10328
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 241704 8984 241756 9036
rect 273444 8984 273496 9036
rect 109316 8916 109368 8968
rect 243544 8916 243596 8968
rect 299020 8916 299072 8968
rect 401324 8916 401376 8968
rect 271236 8236 271288 8288
rect 275284 8236 275336 8288
rect 248788 7624 248840 7676
rect 268384 7624 268436 7676
rect 70308 7556 70360 7608
rect 242164 7556 242216 7608
rect 247592 7556 247644 7608
rect 275100 7556 275152 7608
rect 298100 7556 298152 7608
rect 372896 7556 372948 7608
rect 283104 6876 283156 6928
rect 288992 6876 289044 6928
rect 3424 6808 3476 6860
rect 44824 6808 44876 6860
rect 289084 6808 289136 6860
rect 309048 6808 309100 6860
rect 283012 6740 283064 6792
rect 294880 6740 294932 6792
rect 295524 6740 295576 6792
rect 358728 6740 358780 6792
rect 292488 6672 292540 6724
rect 382372 6672 382424 6724
rect 291016 6604 291068 6656
rect 385960 6604 386012 6656
rect 289268 6536 289320 6588
rect 396540 6536 396592 6588
rect 289636 6468 289688 6520
rect 400128 6468 400180 6520
rect 289452 6400 289504 6452
rect 403624 6400 403676 6452
rect 289360 6332 289412 6384
rect 407212 6332 407264 6384
rect 290924 6264 290976 6316
rect 410800 6264 410852 6316
rect 238116 6196 238168 6248
rect 273352 6196 273404 6248
rect 290740 6196 290792 6248
rect 416688 6196 416740 6248
rect 119896 6128 119948 6180
rect 251640 6128 251692 6180
rect 254676 6128 254728 6180
rect 276480 6128 276532 6180
rect 292396 6128 292448 6180
rect 420184 6128 420236 6180
rect 281816 5516 281868 5568
rect 284208 5516 284260 5568
rect 240508 4904 240560 4956
rect 273260 4904 273312 4956
rect 283472 4904 283524 4956
rect 290188 4904 290240 4956
rect 227536 4836 227588 4888
rect 270500 4836 270552 4888
rect 286324 4836 286376 4888
rect 297272 4836 297324 4888
rect 80888 4768 80940 4820
rect 244556 4768 244608 4820
rect 284300 4768 284352 4820
rect 298468 4768 298520 4820
rect 278320 4156 278372 4208
rect 279424 4156 279476 4208
rect 281724 4156 281776 4208
rect 285404 4156 285456 4208
rect 299572 4156 299624 4208
rect 300768 4156 300820 4208
rect 2872 4088 2924 4140
rect 7564 4088 7616 4140
rect 45468 4088 45520 4140
rect 46296 4088 46348 4140
rect 257068 4088 257120 4140
rect 260196 4088 260248 4140
rect 277124 4088 277176 4140
rect 279516 4088 279568 4140
rect 288348 4088 288400 4140
rect 335084 4088 335136 4140
rect 338764 4088 338816 4140
rect 371700 4088 371752 4140
rect 434444 4088 434496 4140
rect 439136 4088 439188 4140
rect 536196 4088 536248 4140
rect 538404 4088 538456 4140
rect 295340 4020 295392 4072
rect 356336 4020 356388 4072
rect 428464 4020 428516 4072
rect 439412 4020 439464 4072
rect 246396 3952 246448 4004
rect 253296 3952 253348 4004
rect 295432 3952 295484 4004
rect 359924 3952 359976 4004
rect 427268 3952 427320 4004
rect 439228 3952 439280 4004
rect 244096 3884 244148 3936
rect 254584 3884 254636 3936
rect 295248 3884 295300 3936
rect 381176 3884 381228 3936
rect 426164 3884 426216 3936
rect 438860 3884 438912 3936
rect 239312 3816 239364 3868
rect 253388 3816 253440 3868
rect 258172 3816 258224 3868
rect 265624 3816 265676 3868
rect 291108 3816 291160 3868
rect 378876 3816 378928 3868
rect 424968 3816 425020 3868
rect 437664 3816 437716 3868
rect 516784 3816 516836 3868
rect 519544 3816 519596 3868
rect 574744 3816 574796 3868
rect 577412 3816 577464 3868
rect 35992 3748 36044 3800
rect 46204 3748 46256 3800
rect 135260 3748 135312 3800
rect 136456 3748 136508 3800
rect 171968 3748 172020 3800
rect 261392 3748 261444 3800
rect 295156 3748 295208 3800
rect 388260 3748 388312 3800
rect 423772 3748 423824 3800
rect 437848 3748 437900 3800
rect 11152 3680 11204 3732
rect 39304 3680 39356 3732
rect 53748 3680 53800 3732
rect 54484 3680 54536 3732
rect 82084 3680 82136 3732
rect 93124 3680 93176 3732
rect 124680 3680 124732 3732
rect 238024 3680 238076 3732
rect 242900 3680 242952 3732
rect 264244 3680 264296 3732
rect 289728 3680 289780 3732
rect 395344 3680 395396 3732
rect 422576 3680 422628 3732
rect 437480 3680 437532 3732
rect 462964 3680 463016 3732
rect 39580 3612 39632 3664
rect 95884 3612 95936 3664
rect 96252 3612 96304 3664
rect 97264 3612 97316 3664
rect 102232 3612 102284 3664
rect 248696 3612 248748 3664
rect 251180 3612 251232 3664
rect 261484 3612 261536 3664
rect 293500 3612 293552 3664
rect 402520 3612 402572 3664
rect 421380 3612 421432 3664
rect 439044 3612 439096 3664
rect 442264 3612 442316 3664
rect 447416 3612 447468 3664
rect 456064 3612 456116 3664
rect 465172 3612 465224 3664
rect 1676 3544 1728 3596
rect 4804 3544 4856 3596
rect 4068 3476 4120 3528
rect 10324 3544 10376 3596
rect 12348 3544 12400 3596
rect 13084 3544 13136 3596
rect 20628 3544 20680 3596
rect 21364 3544 21416 3596
rect 25320 3544 25372 3596
rect 71044 3544 71096 3596
rect 71504 3544 71556 3596
rect 72424 3544 72476 3596
rect 85672 3544 85724 3596
rect 88984 3544 89036 3596
rect 89260 3544 89312 3596
rect 244740 3544 244792 3596
rect 244832 3544 244884 3596
rect 249984 3544 250036 3596
rect 258172 3544 258224 3596
rect 258264 3544 258316 3596
rect 260104 3544 260156 3596
rect 267740 3544 267792 3596
rect 273904 3544 273956 3596
rect 281448 3544 281500 3596
rect 7656 3476 7708 3528
rect 8944 3476 8996 3528
rect 15936 3476 15988 3528
rect 572 3408 624 3460
rect 25504 3408 25556 3460
rect 27712 3408 27764 3460
rect 31024 3408 31076 3460
rect 33600 3408 33652 3460
rect 35164 3408 35216 3460
rect 38384 3408 38436 3460
rect 39396 3408 39448 3460
rect 40684 3408 40736 3460
rect 43444 3408 43496 3460
rect 46664 3476 46716 3528
rect 47584 3476 47636 3528
rect 47860 3476 47912 3528
rect 48964 3476 49016 3528
rect 56048 3476 56100 3528
rect 57336 3476 57388 3528
rect 60740 3476 60792 3528
rect 61660 3476 61712 3528
rect 83280 3476 83332 3528
rect 253480 3476 253532 3528
rect 269764 3476 269816 3528
rect 281632 3476 281684 3528
rect 283104 3476 283156 3528
rect 293868 3544 293920 3596
rect 406016 3544 406068 3596
rect 418988 3544 419040 3596
rect 438952 3544 439004 3596
rect 443644 3544 443696 3596
rect 292580 3476 292632 3528
rect 295064 3476 295116 3528
rect 409604 3476 409656 3528
rect 417884 3476 417936 3528
rect 437756 3476 437808 3528
rect 440240 3476 440292 3528
rect 441528 3476 441580 3528
rect 448520 3476 448572 3528
rect 449808 3476 449860 3528
rect 453304 3544 453356 3596
rect 455696 3544 455748 3596
rect 467104 3544 467156 3596
rect 469864 3544 469916 3596
rect 480536 3544 480588 3596
rect 471060 3476 471112 3528
rect 471244 3476 471296 3528
rect 473452 3476 473504 3528
rect 476764 3476 476816 3528
rect 484032 3544 484084 3596
rect 491944 3544 491996 3596
rect 494704 3544 494756 3596
rect 500224 3544 500276 3596
rect 501788 3544 501840 3596
rect 511264 3544 511316 3596
rect 513564 3544 513616 3596
rect 514024 3544 514076 3596
rect 515956 3544 516008 3596
rect 549904 3544 549956 3596
rect 551468 3544 551520 3596
rect 481640 3476 481692 3528
rect 482468 3476 482520 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 496084 3476 496136 3528
rect 497096 3476 497148 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 514116 3476 514168 3528
rect 514760 3476 514812 3528
rect 523040 3476 523092 3528
rect 523868 3476 523920 3528
rect 527916 3476 527968 3528
rect 533712 3476 533764 3528
rect 547880 3476 547932 3528
rect 548708 3476 548760 3528
rect 571984 3476 572036 3528
rect 573916 3476 573968 3528
rect 581000 3476 581052 3528
rect 581828 3476 581880 3528
rect 64144 3408 64196 3460
rect 64328 3408 64380 3460
rect 68284 3408 68336 3460
rect 79692 3408 79744 3460
rect 244464 3408 244516 3460
rect 252376 3408 252428 3460
rect 271144 3408 271196 3460
rect 30104 3340 30156 3392
rect 40592 3340 40644 3392
rect 48964 3340 49016 3392
rect 50344 3340 50396 3392
rect 84476 3340 84528 3392
rect 89260 3340 89312 3392
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 262956 3340 263008 3392
rect 269856 3340 269908 3392
rect 292120 3340 292172 3392
rect 413100 3408 413152 3460
rect 415492 3408 415544 3460
rect 437572 3408 437624 3460
rect 450544 3408 450596 3460
rect 452108 3408 452160 3460
rect 456892 3408 456944 3460
rect 458088 3408 458140 3460
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332692 3340 332744 3392
rect 333888 3340 333940 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 430856 3340 430908 3392
rect 438032 3340 438084 3392
rect 445116 3340 445168 3392
rect 569132 3408 569184 3460
rect 570604 3408 570656 3460
rect 572720 3408 572772 3460
rect 57244 3272 57296 3324
rect 58624 3272 58676 3324
rect 65524 3272 65576 3324
rect 66904 3272 66956 3324
rect 259460 3272 259512 3324
rect 264336 3272 264388 3324
rect 435548 3272 435600 3324
rect 439320 3272 439372 3324
rect 6460 3204 6512 3256
rect 7564 3204 7616 3256
rect 78588 3204 78640 3256
rect 82176 3204 82228 3256
rect 478236 3204 478288 3256
rect 479340 3204 479392 3256
rect 554044 3204 554096 3256
rect 557356 3204 557408 3256
rect 293316 3136 293368 3188
rect 296076 3136 296128 3188
rect 433248 3136 433300 3188
rect 440424 3136 440476 3188
rect 485044 3136 485096 3188
rect 487620 3136 487672 3188
rect 534724 3136 534776 3188
rect 537208 3136 537260 3188
rect 560944 3136 560996 3188
rect 563244 3136 563296 3188
rect 567844 3136 567896 3188
rect 570328 3136 570380 3188
rect 19432 3068 19484 3120
rect 22744 3068 22796 3120
rect 273628 3068 273680 3120
rect 278136 3068 278188 3120
rect 270040 3000 270092 3052
rect 272524 3000 272576 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 472624 3000 472676 3052
rect 474556 3000 474608 3052
rect 503076 3000 503128 3052
rect 505376 3000 505428 3052
rect 538864 3000 538916 3052
rect 540796 3000 540848 3052
rect 563704 3000 563756 3052
rect 565636 3000 565688 3052
rect 8760 2932 8812 2984
rect 14464 2932 14516 2984
rect 540244 2932 540296 2984
rect 541992 2932 542044 2984
rect 552756 2932 552808 2984
rect 554964 2932 555016 2984
rect 51356 2864 51408 2916
rect 53104 2864 53156 2916
rect 73804 2864 73856 2916
rect 75184 2864 75236 2916
rect 494796 2864 494848 2916
rect 499396 2864 499448 2916
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3160 553722 3188 553823
rect 3148 553716 3200 553722
rect 3148 553658 3200 553664
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 2870 501800 2926 501809
rect 2870 501735 2926 501744
rect 2884 501022 2912 501735
rect 2872 501016 2924 501022
rect 2872 500958 2924 500964
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 2870 449576 2926 449585
rect 2870 449511 2926 449520
rect 2884 447846 2912 449511
rect 3436 449206 3464 619103
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3528 450634 3556 566879
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3516 450628 3568 450634
rect 3516 450570 3568 450576
rect 3620 450566 3648 514791
rect 4816 467158 4844 683674
rect 6932 471306 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 18604 670744 18656 670750
rect 18604 670686 18656 670692
rect 13084 656940 13136 656946
rect 13084 656882 13136 656888
rect 10324 579692 10376 579698
rect 10324 579634 10376 579640
rect 8944 553716 8996 553722
rect 8944 553658 8996 553664
rect 6920 471300 6972 471306
rect 6920 471242 6972 471248
rect 4804 467152 4856 467158
rect 4804 467094 4856 467100
rect 8956 458862 8984 553658
rect 10336 469878 10364 579634
rect 10324 469872 10376 469878
rect 10324 469814 10376 469820
rect 13096 460222 13124 656882
rect 17224 605872 17276 605878
rect 17224 605814 17276 605820
rect 14464 527196 14516 527202
rect 14464 527138 14516 527144
rect 14476 472666 14504 527138
rect 14464 472660 14516 472666
rect 14464 472602 14516 472608
rect 17236 464370 17264 605814
rect 17224 464364 17276 464370
rect 17224 464306 17276 464312
rect 13084 460216 13136 460222
rect 13084 460158 13136 460164
rect 8944 458856 8996 458862
rect 8944 458798 8996 458804
rect 18616 456074 18644 670686
rect 21364 501016 21416 501022
rect 21364 500958 21416 500964
rect 21376 457502 21404 500958
rect 21364 457496 21416 457502
rect 21364 457438 21416 457444
rect 18604 456068 18656 456074
rect 18604 456010 18656 456016
rect 3608 450560 3660 450566
rect 3608 450502 3660 450508
rect 23492 449274 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 23480 449268 23532 449274
rect 23480 449210 23532 449216
rect 3424 449200 3476 449206
rect 3424 449142 3476 449148
rect 40052 447914 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 478174 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 71780 478168 71832 478174
rect 71780 478110 71832 478116
rect 88352 449410 88380 702406
rect 105464 700330 105492 703520
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 88340 449404 88392 449410
rect 88340 449346 88392 449352
rect 136652 447982 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 153212 449546 153240 702406
rect 166264 700324 166316 700330
rect 166264 700266 166316 700272
rect 166276 468518 166304 700266
rect 166264 468512 166316 468518
rect 166264 468454 166316 468460
rect 169772 465730 169800 702406
rect 198004 632120 198056 632126
rect 198004 632062 198056 632068
rect 198016 474026 198044 632062
rect 198004 474020 198056 474026
rect 198004 473962 198056 473968
rect 169760 465724 169812 465730
rect 169760 465666 169812 465672
rect 153200 449540 153252 449546
rect 153200 449482 153252 449488
rect 201512 448050 201540 702986
rect 217968 700324 218020 700330
rect 217968 700266 218020 700272
rect 217874 516896 217930 516905
rect 217874 516831 217930 516840
rect 217782 515944 217838 515953
rect 217782 515879 217838 515888
rect 217598 513768 217654 513777
rect 217598 513703 217654 513712
rect 217322 488336 217378 488345
rect 217322 488271 217378 488280
rect 217336 478922 217364 488271
rect 217506 488064 217562 488073
rect 217506 487999 217562 488008
rect 217324 478916 217376 478922
rect 217324 478858 217376 478864
rect 217520 476814 217548 487999
rect 217612 478310 217640 513703
rect 217690 489968 217746 489977
rect 217690 489903 217746 489912
rect 217600 478304 217652 478310
rect 217600 478246 217652 478252
rect 217508 476808 217560 476814
rect 217508 476750 217560 476756
rect 217704 451926 217732 489903
rect 217796 472734 217824 515879
rect 217784 472728 217836 472734
rect 217784 472670 217836 472676
rect 217888 471374 217916 516831
rect 217876 471368 217928 471374
rect 217876 471310 217928 471316
rect 217692 451920 217744 451926
rect 217692 451862 217744 451868
rect 201500 448044 201552 448050
rect 201500 447986 201552 447992
rect 136640 447976 136692 447982
rect 136640 447918 136692 447924
rect 40040 447908 40092 447914
rect 40040 447850 40092 447856
rect 2872 447840 2924 447846
rect 2872 447782 2924 447788
rect 57244 446820 57296 446826
rect 57244 446762 57296 446768
rect 7564 444440 7616 444446
rect 7564 444382 7616 444388
rect 3516 443692 3568 443698
rect 3516 443634 3568 443640
rect 3424 423632 3476 423638
rect 3422 423600 3424 423609
rect 3476 423600 3478 423609
rect 3422 423535 3478 423544
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 3424 410576 3476 410582
rect 2962 410544 3018 410553
rect 3424 410518 3476 410524
rect 2962 410479 3018 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3056 372564 3108 372570
rect 3056 372506 3108 372512
rect 3068 371385 3096 372506
rect 3054 371376 3110 371385
rect 3054 371311 3110 371320
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 293956 3384 293962
rect 3332 293898 3384 293904
rect 3344 293185 3372 293898
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 45529 3464 410518
rect 3528 201929 3556 443634
rect 3608 442264 3660 442270
rect 3608 442206 3660 442212
rect 3620 358465 3648 442206
rect 7576 423638 7604 444382
rect 7564 423632 7616 423638
rect 7564 423574 7616 423580
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 44824 309800 44876 309806
rect 44824 309742 44876 309748
rect 31760 308644 31812 308650
rect 31760 308586 31812 308592
rect 27620 308508 27672 308514
rect 27620 308450 27672 308456
rect 23480 308440 23532 308446
rect 23480 308382 23532 308388
rect 7564 304292 7616 304298
rect 7564 304234 7616 304240
rect 4160 262880 4212 262886
rect 4160 262822 4212 262828
rect 3608 246356 3660 246362
rect 3608 246298 3660 246304
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3516 164212 3568 164218
rect 3516 164154 3568 164160
rect 3528 162897 3556 164154
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3620 149841 3648 246298
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 4172 16574 4200 262822
rect 4804 247716 4856 247722
rect 4804 247658 4856 247664
rect 4172 16546 4752 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3538
rect 2884 480 2912 4082
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4724 3482 4752 16546
rect 4816 3602 4844 247658
rect 7576 4146 7604 304234
rect 8944 302932 8996 302938
rect 8944 302874 8996 302880
rect 7656 244928 7708 244934
rect 7656 244870 7708 244876
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 3618 7696 244870
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 7576 3590 7696 3618
rect 4080 480 4108 3470
rect 4724 3454 5304 3482
rect 5276 480 5304 3454
rect 7576 3262 7604 3590
rect 8956 3534 8984 302874
rect 10324 300144 10376 300150
rect 10324 300086 10376 300092
rect 9680 287700 9732 287706
rect 9680 287642 9732 287648
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 6460 3256 6512 3262
rect 6460 3198 6512 3204
rect 7564 3256 7616 3262
rect 7564 3198 7616 3204
rect 6472 480 6500 3198
rect 7668 480 7696 3470
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8772 480 8800 2926
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 287642
rect 10336 3602 10364 300086
rect 13084 289128 13136 289134
rect 13084 289070 13136 289076
rect 12440 249076 12492 249082
rect 12440 249018 12492 249024
rect 12452 16574 12480 249018
rect 12452 16546 13032 16574
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 11164 480 11192 3674
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13004 3482 13032 16546
rect 13096 3602 13124 289070
rect 16580 283620 16632 283626
rect 16580 283562 16632 283568
rect 14464 274032 14516 274038
rect 14464 273974 14516 273980
rect 13820 258732 13872 258738
rect 13820 258674 13872 258680
rect 13832 16574 13860 258674
rect 13832 16546 14320 16574
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13004 3454 13584 3482
rect 13556 480 13584 3454
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 2990 14504 273974
rect 16592 16574 16620 283562
rect 20720 282192 20772 282198
rect 20720 282134 20772 282140
rect 17960 251864 18012 251870
rect 17960 251806 18012 251812
rect 16592 16546 17080 16574
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 15948 480 15976 3470
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 251806
rect 20732 16574 20760 282134
rect 22744 275324 22796 275330
rect 22744 275266 22796 275272
rect 21364 261520 21416 261526
rect 21364 261462 21416 261468
rect 20732 16546 21312 16574
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19444 480 19472 3062
rect 20640 480 20668 3538
rect 21284 3482 21312 16546
rect 21376 3602 21404 261462
rect 22100 250504 22152 250510
rect 22100 250446 22152 250452
rect 22112 16574 22140 250446
rect 22112 16546 22600 16574
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21284 3454 21864 3482
rect 21836 480 21864 3454
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 22756 3126 22784 275266
rect 23492 16574 23520 308382
rect 25504 307080 25556 307086
rect 25504 307022 25556 307028
rect 23492 16546 24256 16574
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 24228 480 24256 16546
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25332 480 25360 3538
rect 25516 3466 25544 307022
rect 26240 280832 26292 280838
rect 26240 280774 26292 280780
rect 25504 3460 25556 3466
rect 25504 3402 25556 3408
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 280774
rect 27632 16574 27660 308450
rect 31024 294636 31076 294642
rect 31024 294578 31076 294584
rect 30380 253224 30432 253230
rect 30380 253166 30432 253172
rect 30392 16574 30420 253166
rect 27632 16546 28488 16574
rect 30392 16546 30880 16574
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 27724 480 27752 3402
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30104 3392 30156 3398
rect 30104 3334 30156 3340
rect 30116 480 30144 3334
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31036 3466 31064 294578
rect 31772 16574 31800 308586
rect 39304 308576 39356 308582
rect 39304 308518 39356 308524
rect 34520 291848 34572 291854
rect 34520 291790 34572 291796
rect 31772 16546 31984 16574
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33612 480 33640 3402
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 291790
rect 35164 278044 35216 278050
rect 35164 277986 35216 277992
rect 35176 3466 35204 277986
rect 35900 276684 35952 276690
rect 35900 276626 35952 276632
rect 35912 16574 35940 276626
rect 35912 16546 36768 16574
rect 35992 3800 36044 3806
rect 35992 3742 36044 3748
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 36004 480 36032 3742
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 39316 3738 39344 308518
rect 43444 301504 43496 301510
rect 43444 301446 43496 301452
rect 41420 290488 41472 290494
rect 41420 290430 41472 290436
rect 39396 284980 39448 284986
rect 39396 284922 39448 284928
rect 39304 3732 39356 3738
rect 39304 3674 39356 3680
rect 39408 3466 39436 284922
rect 40684 279472 40736 279478
rect 40684 279414 40736 279420
rect 40696 6914 40724 279414
rect 41432 16574 41460 290430
rect 42800 260160 42852 260166
rect 42800 260102 42852 260108
rect 41432 16546 41920 16574
rect 40604 6886 40724 6914
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 39396 3460 39448 3466
rect 39396 3402 39448 3408
rect 38396 480 38424 3402
rect 39592 480 39620 3606
rect 40604 3398 40632 6886
rect 40684 3460 40736 3466
rect 40684 3402 40736 3408
rect 40592 3392 40644 3398
rect 40592 3334 40644 3340
rect 40696 480 40724 3402
rect 41892 480 41920 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 260102
rect 43456 3466 43484 301446
rect 44180 275392 44232 275398
rect 44180 275334 44232 275340
rect 44192 16574 44220 275334
rect 44192 16546 44312 16574
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 44284 480 44312 16546
rect 44836 6866 44864 309742
rect 46204 308712 46256 308718
rect 46204 308654 46256 308660
rect 44824 6860 44876 6866
rect 44824 6802 44876 6808
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 45480 480 45508 4082
rect 46216 3806 46244 308654
rect 48964 301572 49016 301578
rect 48964 301514 49016 301520
rect 46296 286340 46348 286346
rect 46296 286282 46348 286288
rect 46308 4146 46336 286282
rect 47584 32428 47636 32434
rect 47584 32370 47636 32376
rect 46296 4140 46348 4146
rect 46296 4082 46348 4088
rect 46204 3800 46256 3806
rect 46204 3742 46256 3748
rect 47596 3534 47624 32370
rect 48976 3534 49004 301514
rect 53104 300212 53156 300218
rect 53104 300154 53156 300160
rect 50344 272536 50396 272542
rect 50344 272478 50396 272484
rect 49700 89004 49752 89010
rect 49700 88946 49752 88952
rect 49712 16574 49740 88946
rect 49712 16546 50200 16574
rect 46664 3528 46716 3534
rect 46664 3470 46716 3476
rect 47584 3528 47636 3534
rect 47584 3470 47636 3476
rect 47860 3528 47912 3534
rect 47860 3470 47912 3476
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 46676 480 46704 3470
rect 47872 480 47900 3470
rect 48964 3392 49016 3398
rect 48964 3334 49016 3340
rect 48976 480 49004 3334
rect 50172 480 50200 16546
rect 50356 3398 50384 272478
rect 52460 271176 52512 271182
rect 52460 271118 52512 271124
rect 52472 16574 52500 271118
rect 52472 16546 52592 16574
rect 50344 3392 50396 3398
rect 50344 3334 50396 3340
rect 51356 2916 51408 2922
rect 51356 2858 51408 2864
rect 51368 480 51396 2858
rect 52564 480 52592 16546
rect 53116 2922 53144 300154
rect 53840 298784 53892 298790
rect 53840 298726 53892 298732
rect 53852 16574 53880 298726
rect 54484 293276 54536 293282
rect 54484 293218 54536 293224
rect 53852 16546 54432 16574
rect 53748 3732 53800 3738
rect 53748 3674 53800 3680
rect 53104 2916 53156 2922
rect 53104 2858 53156 2864
rect 53760 480 53788 3674
rect 54404 3482 54432 16546
rect 54496 3738 54524 293218
rect 57256 97986 57284 446762
rect 217980 446690 218008 700266
rect 218072 478242 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700330 235212 703520
rect 267660 700330 267688 703520
rect 283852 700398 283880 703520
rect 300136 700466 300164 703520
rect 332520 700534 332548 703520
rect 348804 700602 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700596 348844 700602
rect 348792 700538 348844 700544
rect 357624 700596 357676 700602
rect 357624 700538 357676 700544
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 300124 700460 300176 700466
rect 300124 700402 300176 700408
rect 357532 700460 357584 700466
rect 357532 700402 357584 700408
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 357440 700324 357492 700330
rect 357440 700266 357492 700272
rect 219346 512816 219402 512825
rect 219346 512751 219402 512760
rect 219254 511048 219310 511057
rect 219254 510983 219310 510992
rect 219162 509960 219218 509969
rect 219162 509895 219218 509904
rect 219070 508192 219126 508201
rect 219070 508127 219126 508136
rect 218060 478236 218112 478242
rect 218060 478178 218112 478184
rect 219084 475386 219112 508127
rect 219072 475380 219124 475386
rect 219072 475322 219124 475328
rect 219176 474094 219204 509895
rect 219164 474088 219216 474094
rect 219164 474030 219216 474036
rect 219268 461650 219296 510983
rect 219256 461644 219308 461650
rect 219256 461586 219308 461592
rect 219360 454714 219388 512751
rect 220084 478916 220136 478922
rect 220084 478858 220136 478864
rect 219348 454708 219400 454714
rect 219348 454650 219400 454656
rect 217968 446684 218020 446690
rect 217968 446626 218020 446632
rect 220096 446486 220124 478858
rect 248420 478304 248472 478310
rect 248420 478246 248472 478252
rect 309140 478304 309192 478310
rect 309140 478246 309192 478252
rect 242898 476912 242954 476921
rect 242898 476847 242954 476856
rect 247038 476912 247094 476921
rect 247038 476847 247094 476856
rect 230480 476808 230532 476814
rect 238852 476808 238904 476814
rect 230480 476750 230532 476756
rect 238758 476776 238814 476785
rect 230492 460934 230520 476750
rect 237472 476740 237524 476746
rect 238852 476750 238904 476756
rect 238758 476711 238760 476720
rect 237472 476682 237524 476688
rect 238812 476711 238814 476720
rect 238760 476682 238812 476688
rect 233240 476672 233292 476678
rect 233240 476614 233292 476620
rect 231860 476332 231912 476338
rect 231860 476274 231912 476280
rect 230492 460906 230704 460934
rect 220084 446480 220136 446486
rect 220084 446422 220136 446428
rect 230388 446480 230440 446486
rect 230388 446422 230440 446428
rect 229836 446072 229888 446078
rect 229836 446014 229888 446020
rect 228364 446004 228416 446010
rect 228364 445946 228416 445952
rect 225696 445188 225748 445194
rect 225696 445130 225748 445136
rect 224224 444984 224276 444990
rect 224224 444926 224276 444932
rect 86224 444712 86276 444718
rect 86224 444654 86276 444660
rect 84844 444644 84896 444650
rect 84844 444586 84896 444592
rect 82084 444576 82136 444582
rect 82084 444518 82136 444524
rect 80704 444508 80756 444514
rect 80704 444450 80756 444456
rect 79324 443012 79376 443018
rect 79324 442954 79376 442960
rect 71044 308848 71096 308854
rect 71044 308790 71096 308796
rect 64144 308780 64196 308786
rect 64144 308722 64196 308728
rect 57980 307148 58032 307154
rect 57980 307090 58032 307096
rect 57336 269816 57388 269822
rect 57336 269758 57388 269764
rect 57244 97980 57296 97986
rect 57244 97922 57296 97928
rect 54484 3732 54536 3738
rect 54484 3674 54536 3680
rect 57348 3534 57376 269758
rect 57992 16574 58020 307090
rect 60740 297424 60792 297430
rect 60740 297366 60792 297372
rect 58624 289196 58676 289202
rect 58624 289138 58676 289144
rect 57992 16546 58480 16574
rect 56048 3528 56100 3534
rect 54404 3454 54984 3482
rect 56048 3470 56100 3476
rect 57336 3528 57388 3534
rect 57336 3470 57388 3476
rect 54956 480 54984 3454
rect 56060 480 56088 3470
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57256 480 57284 3266
rect 58452 480 58480 16546
rect 58636 3330 58664 289138
rect 59360 268388 59412 268394
rect 59360 268330 59412 268336
rect 58624 3324 58676 3330
rect 58624 3266 58676 3272
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59372 354 59400 268330
rect 60752 3534 60780 297366
rect 62120 265668 62172 265674
rect 62120 265610 62172 265616
rect 62132 16574 62160 265610
rect 62132 16546 63264 16574
rect 60832 10328 60884 10334
rect 60832 10270 60884 10276
rect 60740 3528 60792 3534
rect 60740 3470 60792 3476
rect 60844 480 60872 10270
rect 61660 3528 61712 3534
rect 61660 3470 61712 3476
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3470
rect 63236 480 63264 16546
rect 64156 3466 64184 308722
rect 68284 307216 68336 307222
rect 68284 307158 68336 307164
rect 66904 295996 66956 296002
rect 66904 295938 66956 295944
rect 66260 264240 66312 264246
rect 66260 264182 66312 264188
rect 66272 16574 66300 264182
rect 66272 16546 66760 16574
rect 64144 3460 64196 3466
rect 64144 3402 64196 3408
rect 64328 3460 64380 3466
rect 64328 3402 64380 3408
rect 64340 480 64368 3402
rect 65524 3324 65576 3330
rect 65524 3266 65576 3272
rect 65536 480 65564 3266
rect 66732 480 66760 16546
rect 66916 3330 66944 295938
rect 67640 283688 67692 283694
rect 67640 283630 67692 283636
rect 66904 3324 66956 3330
rect 66904 3266 66956 3272
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 283630
rect 68296 3466 68324 307158
rect 69020 294704 69072 294710
rect 69020 294646 69072 294652
rect 69032 16574 69060 294646
rect 69032 16546 69152 16574
rect 68284 3460 68336 3466
rect 68284 3402 68336 3408
rect 69124 480 69152 16546
rect 70308 7608 70360 7614
rect 70308 7550 70360 7556
rect 70320 480 70348 7550
rect 71056 3602 71084 308790
rect 75920 305720 75972 305726
rect 75920 305662 75972 305668
rect 72424 305652 72476 305658
rect 72424 305594 72476 305600
rect 71780 291916 71832 291922
rect 71780 291858 71832 291864
rect 71792 16574 71820 291858
rect 71792 16546 72372 16574
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 71504 3596 71556 3602
rect 71504 3538 71556 3544
rect 71516 480 71544 3538
rect 72344 3482 72372 16546
rect 72436 3602 72464 305594
rect 74540 282260 74592 282266
rect 74540 282202 74592 282208
rect 74552 16574 74580 282202
rect 75184 262948 75236 262954
rect 75184 262890 75236 262896
rect 74552 16546 75040 16574
rect 72424 3596 72476 3602
rect 72424 3538 72476 3544
rect 72344 3454 72648 3482
rect 72620 480 72648 3454
rect 73804 2916 73856 2922
rect 73804 2858 73856 2864
rect 73816 480 73844 2858
rect 75012 480 75040 16546
rect 75196 2922 75224 262890
rect 75184 2916 75236 2922
rect 75184 2858 75236 2864
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 305662
rect 77300 261588 77352 261594
rect 77300 261530 77352 261536
rect 77312 16574 77340 261530
rect 79336 85542 79364 442954
rect 80716 137970 80744 444450
rect 80704 137964 80756 137970
rect 80704 137906 80756 137912
rect 82096 111790 82124 444518
rect 82176 304360 82228 304366
rect 82176 304302 82228 304308
rect 82084 111784 82136 111790
rect 82084 111726 82136 111732
rect 79324 85536 79376 85542
rect 79324 85478 79376 85484
rect 77312 16546 77432 16574
rect 77404 480 77432 16546
rect 80888 4820 80940 4826
rect 80888 4762 80940 4768
rect 79692 3460 79744 3466
rect 79692 3402 79744 3408
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 78600 480 78628 3198
rect 79704 480 79732 3402
rect 80900 480 80928 4762
rect 82084 3732 82136 3738
rect 82084 3674 82136 3680
rect 82096 480 82124 3674
rect 82188 3262 82216 304302
rect 84856 164218 84884 444586
rect 85580 304428 85632 304434
rect 85580 304370 85632 304376
rect 84844 164212 84896 164218
rect 84844 164154 84896 164160
rect 85592 16574 85620 304370
rect 86236 215286 86264 444654
rect 220084 443420 220136 443426
rect 220084 443362 220136 443368
rect 98644 443148 98696 443154
rect 98644 443090 98696 443096
rect 95976 443080 96028 443086
rect 95976 443022 96028 443028
rect 95884 308984 95936 308990
rect 95884 308926 95936 308932
rect 93124 303068 93176 303074
rect 93124 303010 93176 303016
rect 86960 297492 87012 297498
rect 86960 297434 87012 297440
rect 86224 215280 86276 215286
rect 86224 215222 86276 215228
rect 86972 16574 87000 297434
rect 89720 286408 89772 286414
rect 89720 286350 89772 286356
rect 88984 280900 89036 280906
rect 88984 280842 89036 280848
rect 88340 254584 88392 254590
rect 88340 254526 88392 254532
rect 88352 16574 88380 254526
rect 85592 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 88932 16574
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 82176 3256 82228 3262
rect 82176 3198 82228 3204
rect 83292 480 83320 3470
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 84488 480 84516 3334
rect 85684 480 85712 3538
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 88904 3482 88932 16546
rect 88996 3602 89024 280842
rect 89732 16574 89760 286350
rect 92480 279540 92532 279546
rect 92480 279482 92532 279488
rect 91100 258800 91152 258806
rect 91100 258742 91152 258748
rect 91112 16574 91140 258742
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 88984 3596 89036 3602
rect 88984 3538 89036 3544
rect 89260 3596 89312 3602
rect 89260 3538 89312 3544
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 89272 3398 89300 3538
rect 89260 3392 89312 3398
rect 89260 3334 89312 3340
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 279482
rect 93136 3738 93164 303010
rect 93860 303000 93912 303006
rect 93860 302942 93912 302948
rect 93872 6914 93900 302942
rect 93952 296064 94004 296070
rect 93952 296006 94004 296012
rect 93964 16574 93992 296006
rect 93964 16546 94728 16574
rect 93872 6886 93992 6914
rect 93124 3732 93176 3738
rect 93124 3674 93176 3680
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95896 3670 95924 308926
rect 95988 189038 96016 443022
rect 97264 308916 97316 308922
rect 97264 308858 97316 308864
rect 96620 285048 96672 285054
rect 96620 284990 96672 284996
rect 95976 189032 96028 189038
rect 95976 188974 96028 188980
rect 96632 16574 96660 284990
rect 96632 16546 97212 16574
rect 95884 3664 95936 3670
rect 95884 3606 95936 3612
rect 96252 3664 96304 3670
rect 96252 3606 96304 3612
rect 96264 480 96292 3606
rect 97184 3482 97212 16546
rect 97276 3670 97304 308858
rect 98000 253292 98052 253298
rect 98000 253234 98052 253240
rect 97816 243568 97868 243574
rect 97816 243510 97868 243516
rect 97724 243432 97776 243438
rect 97724 243374 97776 243380
rect 97736 196897 97764 243374
rect 97722 196888 97778 196897
rect 97722 196823 97778 196832
rect 97828 195945 97856 243510
rect 97908 243500 97960 243506
rect 97908 243442 97960 243448
rect 97814 195936 97870 195945
rect 97814 195871 97870 195880
rect 97814 193760 97870 193769
rect 97814 193695 97870 193704
rect 97538 192808 97594 192817
rect 97538 192743 97594 192752
rect 97446 168328 97502 168337
rect 97446 168263 97502 168272
rect 97460 159730 97488 168263
rect 97552 159798 97580 192743
rect 97630 191040 97686 191049
rect 97630 190975 97686 190984
rect 97644 159866 97672 190975
rect 97722 189952 97778 189961
rect 97722 189887 97778 189896
rect 97632 159860 97684 159866
rect 97632 159802 97684 159808
rect 97540 159792 97592 159798
rect 97540 159734 97592 159740
rect 97448 159724 97500 159730
rect 97448 159666 97500 159672
rect 97736 157690 97764 189887
rect 97828 159934 97856 193695
rect 97920 188193 97948 243442
rect 97906 188184 97962 188193
rect 97906 188119 97962 188128
rect 97906 169960 97962 169969
rect 97906 169895 97962 169904
rect 97816 159928 97868 159934
rect 97816 159870 97868 159876
rect 97920 159662 97948 169895
rect 97908 159656 97960 159662
rect 97908 159598 97960 159604
rect 97724 157684 97776 157690
rect 97724 157626 97776 157632
rect 98012 16574 98040 253234
rect 98656 241466 98684 443090
rect 99288 273964 99340 273970
rect 99288 273906 99340 273912
rect 98644 241460 98696 241466
rect 98644 241402 98696 241408
rect 99300 168065 99328 273906
rect 220096 255270 220124 443362
rect 221464 443284 221516 443290
rect 221464 443226 221516 443232
rect 221476 346390 221504 443226
rect 221464 346384 221516 346390
rect 221464 346326 221516 346332
rect 224236 267714 224264 444926
rect 225604 443488 225656 443494
rect 225604 443430 225656 443436
rect 225616 306338 225644 443430
rect 225708 320142 225736 445130
rect 226984 443556 227036 443562
rect 226984 443498 227036 443504
rect 226996 411262 227024 443498
rect 226984 411256 227036 411262
rect 226984 411198 227036 411204
rect 225696 320136 225748 320142
rect 225696 320078 225748 320084
rect 225604 306332 225656 306338
rect 225604 306274 225656 306280
rect 224224 267708 224276 267714
rect 224224 267650 224276 267656
rect 220084 255264 220136 255270
rect 220084 255206 220136 255212
rect 228376 246362 228404 445946
rect 229744 445936 229796 445942
rect 229744 445878 229796 445884
rect 228548 445256 228600 445262
rect 228548 445198 228600 445204
rect 228456 444916 228508 444922
rect 228456 444858 228508 444864
rect 228468 293962 228496 444858
rect 228560 372570 228588 445198
rect 228640 443352 228692 443358
rect 228640 443294 228692 443300
rect 228652 398818 228680 443294
rect 229756 410582 229784 445878
rect 229848 442270 229876 446014
rect 230400 443564 230428 446422
rect 230676 443578 230704 460906
rect 231872 447098 231900 476274
rect 231952 451920 232004 451926
rect 231952 451862 232004 451868
rect 231860 447092 231912 447098
rect 231860 447034 231912 447040
rect 231964 443578 231992 451862
rect 232412 447092 232464 447098
rect 232412 447034 232464 447040
rect 230676 443550 231150 443578
rect 231886 443550 231992 443578
rect 232424 443578 232452 447034
rect 233252 443578 233280 476614
rect 233332 476604 233384 476610
rect 233332 476546 233384 476552
rect 233344 460934 233372 476546
rect 235920 476474 236040 476490
rect 235920 476468 236052 476474
rect 235920 476462 236000 476468
rect 234620 476196 234672 476202
rect 234620 476138 234672 476144
rect 233344 460906 233832 460934
rect 233804 443578 233832 460906
rect 234632 443578 234660 476138
rect 234712 476128 234764 476134
rect 234712 476070 234764 476076
rect 234724 460934 234752 476070
rect 235920 475946 235948 476462
rect 236000 476410 236052 476416
rect 235998 476368 236054 476377
rect 235998 476303 236000 476312
rect 236052 476303 236054 476312
rect 236092 476332 236144 476338
rect 236000 476274 236052 476280
rect 236092 476274 236144 476280
rect 235998 476232 236054 476241
rect 235998 476167 236054 476176
rect 236012 476134 236040 476167
rect 236000 476128 236052 476134
rect 236000 476070 236052 476076
rect 235920 475918 236040 475946
rect 234724 460906 235488 460934
rect 235460 443578 235488 460906
rect 236012 447098 236040 475918
rect 236104 460934 236132 476274
rect 237378 476232 237434 476241
rect 237378 476167 237380 476176
rect 237432 476167 237434 476176
rect 237380 476138 237432 476144
rect 237484 470594 237512 476682
rect 238864 476610 238892 476750
rect 242912 476746 242940 476847
rect 247052 476814 247080 476847
rect 247040 476808 247092 476814
rect 247040 476750 247092 476756
rect 242900 476740 242952 476746
rect 242900 476682 242952 476688
rect 238852 476604 238904 476610
rect 238852 476546 238904 476552
rect 242900 476536 242952 476542
rect 245752 476536 245804 476542
rect 242900 476478 242952 476484
rect 244370 476504 244426 476513
rect 240140 476468 240192 476474
rect 240140 476410 240192 476416
rect 238944 476264 238996 476270
rect 238944 476206 238996 476212
rect 238852 475380 238904 475386
rect 238852 475322 238904 475328
rect 237392 470566 237512 470594
rect 237392 460934 237420 470566
rect 236104 460906 236224 460934
rect 237392 460906 237696 460934
rect 236000 447092 236052 447098
rect 236000 447034 236052 447040
rect 236196 443578 236224 460906
rect 237012 447092 237064 447098
rect 237012 447034 237064 447040
rect 237024 443578 237052 447034
rect 237668 443578 237696 460906
rect 232424 443550 232714 443578
rect 233252 443550 233450 443578
rect 233804 443550 234278 443578
rect 234632 443550 235014 443578
rect 235460 443550 235842 443578
rect 236196 443550 236578 443578
rect 237024 443550 237314 443578
rect 237668 443550 238142 443578
rect 238864 443564 238892 475322
rect 238956 460934 238984 476206
rect 238956 460906 239352 460934
rect 239324 443578 239352 460906
rect 240152 443578 240180 476410
rect 240230 476232 240286 476241
rect 242806 476232 242862 476241
rect 240230 476167 240286 476176
rect 241520 476196 241572 476202
rect 240244 460934 240272 476167
rect 242806 476167 242862 476176
rect 241520 476138 241572 476144
rect 240244 460906 240824 460934
rect 240796 443578 240824 460906
rect 241532 447098 241560 476138
rect 242820 476134 242848 476167
rect 242808 476128 242860 476134
rect 242808 476070 242860 476076
rect 241612 474088 241664 474094
rect 241612 474030 241664 474036
rect 241520 447092 241572 447098
rect 241520 447034 241572 447040
rect 241624 443578 241652 474030
rect 242912 460934 242940 476478
rect 248432 476490 248460 478246
rect 249798 477320 249854 477329
rect 249798 477255 249854 477264
rect 268014 477320 268070 477329
rect 268014 477255 268070 477264
rect 249812 476678 249840 477255
rect 258078 477048 258134 477057
rect 258078 476983 258134 476992
rect 252742 476912 252798 476921
rect 252742 476847 252798 476856
rect 255410 476912 255466 476921
rect 255410 476847 255466 476856
rect 249800 476672 249852 476678
rect 249800 476614 249852 476620
rect 251180 476672 251232 476678
rect 251180 476614 251232 476620
rect 248604 476604 248656 476610
rect 248604 476546 248656 476552
rect 245752 476478 245804 476484
rect 244370 476439 244426 476448
rect 244278 476368 244334 476377
rect 244278 476303 244280 476312
rect 244332 476303 244334 476312
rect 244280 476274 244332 476280
rect 244384 476270 244412 476439
rect 244372 476264 244424 476270
rect 244372 476206 244424 476212
rect 245658 476232 245714 476241
rect 245658 476167 245660 476176
rect 245712 476167 245714 476176
rect 245660 476138 245712 476144
rect 244280 476128 244332 476134
rect 244280 476070 244332 476076
rect 242912 460906 243216 460934
rect 242348 447092 242400 447098
rect 242348 447034 242400 447040
rect 242360 443578 242388 447034
rect 243188 443578 243216 460906
rect 239324 443550 239706 443578
rect 240152 443550 240442 443578
rect 240796 443550 241270 443578
rect 241624 443550 242006 443578
rect 242360 443550 242742 443578
rect 243188 443550 243570 443578
rect 244292 443564 244320 476070
rect 244372 461644 244424 461650
rect 244372 461586 244424 461592
rect 244384 460934 244412 461586
rect 244384 460906 244688 460934
rect 244372 446140 244424 446146
rect 244372 446082 244424 446088
rect 244384 443698 244412 446082
rect 244372 443692 244424 443698
rect 244372 443634 244424 443640
rect 244660 443578 244688 460906
rect 245764 447098 245792 476478
rect 248340 476462 248460 476490
rect 247316 476332 247368 476338
rect 247316 476274 247368 476280
rect 247038 476232 247094 476241
rect 247038 476167 247094 476176
rect 247052 476134 247080 476167
rect 245844 476128 245896 476134
rect 245844 476070 245896 476076
rect 247040 476128 247092 476134
rect 247040 476070 247092 476076
rect 245752 447092 245804 447098
rect 245752 447034 245804 447040
rect 244660 443550 245134 443578
rect 245856 443564 245884 476070
rect 247328 460934 247356 476274
rect 248340 476218 248368 476462
rect 248510 476368 248566 476377
rect 248510 476303 248512 476312
rect 248564 476303 248566 476312
rect 248512 476274 248564 476280
rect 248340 476190 248460 476218
rect 247328 460906 247816 460934
rect 247132 454708 247184 454714
rect 247132 454650 247184 454656
rect 246396 447092 246448 447098
rect 246396 447034 246448 447040
rect 246408 443578 246436 447034
rect 247144 443578 247172 454650
rect 247788 443578 247816 460906
rect 248432 447098 248460 476190
rect 248616 470594 248644 476546
rect 249890 476232 249946 476241
rect 249890 476167 249946 476176
rect 248524 470566 248644 470594
rect 248420 447092 248472 447098
rect 248420 447034 248472 447040
rect 248524 443578 248552 470566
rect 249904 460934 249932 476167
rect 249904 460906 250208 460934
rect 249340 447092 249392 447098
rect 249340 447034 249392 447040
rect 249352 443578 249380 447034
rect 250180 443578 250208 460906
rect 251192 443578 251220 476614
rect 252560 476400 252612 476406
rect 252466 476368 252522 476377
rect 252560 476342 252612 476348
rect 252466 476303 252522 476312
rect 252480 476134 252508 476303
rect 252468 476128 252520 476134
rect 252468 476070 252520 476076
rect 251272 472728 251324 472734
rect 251272 472670 251324 472676
rect 251284 460934 251312 472670
rect 251284 460906 251680 460934
rect 251652 443578 251680 460906
rect 252572 447098 252600 476342
rect 252756 476270 252784 476847
rect 255320 476468 255372 476474
rect 255320 476410 255372 476416
rect 252744 476264 252796 476270
rect 252650 476232 252706 476241
rect 252744 476206 252796 476212
rect 253846 476232 253902 476241
rect 252650 476167 252706 476176
rect 253846 476167 253848 476176
rect 252560 447092 252612 447098
rect 252560 447034 252612 447040
rect 252664 443578 252692 476167
rect 253900 476167 253902 476176
rect 253848 476138 253900 476144
rect 253940 476128 253992 476134
rect 253940 476070 253992 476076
rect 253204 447092 253256 447098
rect 253204 447034 253256 447040
rect 253216 443578 253244 447034
rect 253952 445466 253980 476070
rect 254032 471368 254084 471374
rect 254032 471310 254084 471316
rect 253940 445460 253992 445466
rect 253940 445402 253992 445408
rect 254044 443578 254072 471310
rect 255332 460934 255360 476410
rect 255424 476338 255452 476847
rect 255962 476368 256018 476377
rect 255412 476332 255464 476338
rect 255962 476303 256018 476312
rect 256792 476332 256844 476338
rect 255412 476274 255464 476280
rect 255332 460906 255544 460934
rect 254860 445460 254912 445466
rect 254860 445402 254912 445408
rect 254872 443578 254900 445402
rect 255516 443578 255544 460906
rect 255976 447098 256004 476303
rect 256792 476274 256844 476280
rect 256606 476232 256662 476241
rect 256606 476167 256662 476176
rect 256700 476196 256752 476202
rect 255964 447092 256016 447098
rect 255964 447034 256016 447040
rect 256620 447030 256648 476167
rect 256700 476138 256752 476144
rect 256608 447024 256660 447030
rect 256608 446966 256660 446972
rect 246408 443550 246698 443578
rect 247144 443550 247434 443578
rect 247788 443550 248170 443578
rect 248524 443550 248998 443578
rect 249352 443550 249734 443578
rect 250180 443550 250562 443578
rect 251192 443550 251298 443578
rect 251652 443550 252126 443578
rect 252664 443550 252862 443578
rect 253216 443550 253598 443578
rect 254044 443550 254426 443578
rect 254872 443550 255162 443578
rect 255516 443550 255990 443578
rect 256712 443564 256740 476138
rect 256804 460934 256832 476274
rect 258092 476134 258120 476983
rect 258722 476776 258778 476785
rect 258722 476711 258778 476720
rect 263598 476776 263654 476785
rect 263598 476711 263654 476720
rect 258262 476640 258318 476649
rect 258262 476575 258318 476584
rect 258276 476542 258304 476575
rect 258264 476536 258316 476542
rect 258264 476478 258316 476484
rect 258172 476264 258224 476270
rect 258172 476206 258224 476212
rect 258080 476128 258132 476134
rect 258080 476070 258132 476076
rect 258184 460934 258212 476206
rect 256804 460906 257200 460934
rect 258184 460906 258672 460934
rect 257172 443578 257200 460906
rect 258264 447092 258316 447098
rect 258264 447034 258316 447040
rect 257172 443550 257554 443578
rect 258276 443564 258304 447034
rect 258644 443578 258672 460906
rect 258736 447098 258764 476711
rect 263612 476678 263640 476711
rect 263600 476672 263652 476678
rect 260838 476640 260894 476649
rect 263600 476614 263652 476620
rect 260838 476575 260840 476584
rect 260892 476575 260894 476584
rect 260840 476546 260892 476552
rect 259552 476536 259604 476542
rect 259552 476478 259604 476484
rect 264242 476504 264298 476513
rect 259564 460934 259592 476478
rect 264242 476439 264298 476448
rect 264978 476504 265034 476513
rect 268028 476474 268056 477255
rect 270498 477048 270554 477057
rect 270498 476983 270554 476992
rect 304998 477048 305054 477057
rect 304998 476983 305054 476992
rect 307758 477048 307814 477057
rect 307758 476983 307814 476992
rect 264978 476439 265034 476448
rect 268016 476468 268068 476474
rect 261482 476368 261538 476377
rect 261482 476303 261538 476312
rect 260746 476232 260802 476241
rect 260746 476167 260802 476176
rect 260932 476196 260984 476202
rect 259564 460906 260144 460934
rect 258724 447092 258776 447098
rect 258724 447034 258776 447040
rect 259828 447024 259880 447030
rect 259828 446966 259880 446972
rect 258644 443550 259026 443578
rect 259840 443564 259868 446966
rect 260116 443578 260144 460906
rect 260760 447030 260788 476167
rect 260932 476138 260984 476144
rect 260944 460934 260972 476138
rect 260944 460906 261432 460934
rect 261116 447092 261168 447098
rect 261116 447034 261168 447040
rect 260748 447024 260800 447030
rect 260748 446966 260800 446972
rect 261128 443578 261156 447034
rect 261404 445482 261432 460906
rect 261496 446554 261524 476303
rect 262862 476232 262918 476241
rect 262862 476167 262918 476176
rect 262220 476128 262272 476134
rect 262220 476070 262272 476076
rect 262232 460934 262260 476070
rect 262232 460906 262536 460934
rect 261484 446548 261536 446554
rect 261484 446490 261536 446496
rect 261404 445454 261800 445482
rect 261772 443578 261800 445454
rect 262508 443578 262536 460906
rect 262876 447098 262904 476167
rect 263692 461644 263744 461650
rect 263692 461586 263744 461592
rect 262864 447092 262916 447098
rect 262864 447034 262916 447040
rect 260116 443550 260590 443578
rect 261128 443550 261418 443578
rect 261772 443550 262154 443578
rect 262508 443550 262982 443578
rect 263704 443564 263732 461586
rect 264256 446962 264284 476439
rect 264992 476406 265020 476439
rect 268016 476410 268068 476416
rect 264980 476400 265032 476406
rect 264980 476342 265032 476348
rect 265622 476368 265678 476377
rect 265622 476303 265678 476312
rect 267554 476368 267610 476377
rect 270512 476338 270540 476983
rect 277950 476912 278006 476921
rect 277950 476847 278006 476856
rect 302238 476912 302294 476921
rect 302238 476847 302294 476856
rect 276018 476640 276074 476649
rect 276018 476575 276074 476584
rect 276032 476542 276060 476575
rect 276020 476536 276072 476542
rect 276020 476478 276072 476484
rect 273258 476368 273314 476377
rect 267554 476303 267610 476312
rect 270500 476332 270552 476338
rect 265072 456136 265124 456142
rect 265072 456078 265124 456084
rect 264520 447024 264572 447030
rect 264520 446966 264572 446972
rect 264244 446956 264296 446962
rect 264244 446898 264296 446904
rect 264532 443564 264560 446966
rect 265084 443578 265112 456078
rect 265636 446486 265664 476303
rect 266266 476232 266322 476241
rect 266266 476167 266322 476176
rect 266280 451994 266308 476167
rect 267568 475386 267596 476303
rect 273258 476303 273314 476312
rect 274454 476368 274510 476377
rect 274454 476303 274510 476312
rect 270500 476274 270552 476280
rect 273272 476270 273300 476303
rect 273260 476264 273312 476270
rect 267646 476232 267702 476241
rect 267646 476167 267702 476176
rect 269026 476232 269082 476241
rect 269026 476167 269082 476176
rect 270406 476232 270462 476241
rect 270406 476167 270462 476176
rect 271786 476232 271842 476241
rect 271786 476167 271842 476176
rect 273166 476232 273222 476241
rect 273260 476206 273312 476212
rect 273166 476167 273222 476176
rect 267556 475380 267608 475386
rect 267556 475322 267608 475328
rect 266452 463004 266504 463010
rect 266452 462946 266504 462952
rect 266268 451988 266320 451994
rect 266268 451930 266320 451936
rect 265992 446548 266044 446554
rect 265992 446490 266044 446496
rect 265624 446480 265676 446486
rect 265624 446422 265676 446428
rect 265084 443550 265282 443578
rect 266004 443564 266032 446490
rect 266464 443578 266492 462946
rect 267660 453422 267688 476167
rect 268016 457564 268068 457570
rect 268016 457506 268068 457512
rect 267648 453416 267700 453422
rect 267648 453358 267700 453364
rect 267556 447092 267608 447098
rect 267556 447034 267608 447040
rect 266464 443550 266846 443578
rect 267568 443564 267596 447034
rect 268028 443578 268056 457506
rect 269040 455394 269068 476167
rect 269488 458924 269540 458930
rect 269488 458866 269540 458872
rect 269028 455388 269080 455394
rect 269028 455330 269080 455336
rect 269120 446956 269172 446962
rect 269120 446898 269172 446904
rect 268028 443550 268410 443578
rect 269132 443564 269160 446898
rect 269500 443578 269528 458866
rect 270420 451926 270448 476167
rect 270960 453348 271012 453354
rect 270960 453290 271012 453296
rect 270408 451920 270460 451926
rect 270408 451862 270460 451868
rect 270684 446480 270736 446486
rect 270684 446422 270736 446428
rect 269500 443550 269974 443578
rect 270696 443564 270724 446422
rect 270972 443578 271000 453290
rect 271800 452810 271828 476167
rect 271880 460284 271932 460290
rect 271880 460226 271932 460232
rect 271788 452804 271840 452810
rect 271788 452746 271840 452752
rect 271892 447098 271920 460226
rect 273180 451994 273208 476167
rect 274468 474094 274496 476303
rect 274546 476232 274602 476241
rect 274546 476167 274602 476176
rect 275926 476232 275982 476241
rect 275926 476167 275982 476176
rect 277306 476232 277362 476241
rect 277964 476202 277992 476847
rect 291200 476740 291252 476746
rect 291200 476682 291252 476688
rect 278780 476672 278832 476678
rect 278780 476614 278832 476620
rect 278686 476232 278742 476241
rect 277306 476167 277362 476176
rect 277952 476196 278004 476202
rect 274456 474088 274508 474094
rect 274456 474030 274508 474036
rect 273260 464432 273312 464438
rect 273260 464374 273312 464380
rect 271972 451988 272024 451994
rect 271972 451930 272024 451936
rect 273168 451988 273220 451994
rect 273168 451930 273220 451936
rect 271880 447092 271932 447098
rect 271880 447034 271932 447040
rect 271984 443578 272012 451930
rect 273272 447098 273300 464374
rect 274560 454782 274588 476167
rect 274640 475380 274692 475386
rect 274640 475322 274692 475328
rect 274652 460934 274680 475322
rect 275940 461718 275968 476167
rect 276020 465792 276072 465798
rect 276020 465734 276072 465740
rect 275928 461712 275980 461718
rect 275928 461654 275980 461660
rect 274652 460906 275048 460934
rect 274548 454776 274600 454782
rect 274548 454718 274600 454724
rect 273352 453416 273404 453422
rect 273352 453358 273404 453364
rect 272708 447092 272760 447098
rect 272708 447034 272760 447040
rect 273260 447092 273312 447098
rect 273260 447034 273312 447040
rect 272720 443578 272748 447034
rect 273364 443578 273392 453358
rect 274180 447092 274232 447098
rect 274180 447034 274232 447040
rect 274192 443578 274220 447034
rect 275020 443578 275048 460906
rect 276032 443578 276060 465734
rect 276480 455388 276532 455394
rect 276480 455330 276532 455336
rect 276492 443578 276520 455330
rect 277320 453422 277348 476167
rect 278686 476167 278742 476176
rect 277952 476138 278004 476144
rect 277584 476128 277636 476134
rect 277584 476070 277636 476076
rect 277308 453416 277360 453422
rect 277308 453358 277360 453364
rect 277492 451920 277544 451926
rect 277492 451862 277544 451868
rect 277504 447098 277532 451862
rect 277492 447092 277544 447098
rect 277492 447034 277544 447040
rect 277596 443578 277624 476070
rect 278700 451926 278728 476167
rect 278688 451920 278740 451926
rect 278688 451862 278740 451868
rect 278044 447092 278096 447098
rect 278044 447034 278096 447040
rect 278056 443578 278084 447034
rect 278792 443578 278820 476614
rect 280160 476604 280212 476610
rect 280160 476546 280212 476552
rect 280066 476232 280122 476241
rect 280066 476167 280122 476176
rect 280080 454714 280108 476167
rect 280172 460934 280200 476546
rect 281540 476536 281592 476542
rect 281540 476478 281592 476484
rect 280250 476232 280306 476241
rect 280250 476167 280306 476176
rect 280264 461650 280292 476167
rect 280252 461644 280304 461650
rect 280252 461586 280304 461592
rect 280172 460906 280384 460934
rect 280068 454708 280120 454714
rect 280068 454650 280120 454656
rect 279608 452804 279660 452810
rect 279608 452746 279660 452752
rect 279620 443578 279648 452746
rect 280356 443578 280384 460906
rect 281552 447098 281580 476478
rect 282920 476468 282972 476474
rect 282920 476410 282972 476416
rect 281724 451988 281776 451994
rect 281724 451930 281776 451936
rect 281540 447092 281592 447098
rect 281540 447034 281592 447040
rect 281736 443578 281764 451930
rect 282932 447098 282960 476410
rect 284300 476400 284352 476406
rect 284300 476342 284352 476348
rect 283010 476232 283066 476241
rect 283010 476167 283066 476176
rect 283024 456142 283052 476167
rect 283012 456136 283064 456142
rect 283012 456078 283064 456084
rect 283012 454776 283064 454782
rect 283012 454718 283064 454724
rect 281908 447092 281960 447098
rect 281908 447034 281960 447040
rect 282920 447092 282972 447098
rect 282920 447034 282972 447040
rect 270972 443550 271446 443578
rect 271984 443550 272274 443578
rect 272720 443550 273010 443578
rect 273364 443550 273838 443578
rect 274192 443550 274574 443578
rect 275020 443550 275402 443578
rect 276032 443550 276138 443578
rect 276492 443550 276874 443578
rect 277596 443550 277702 443578
rect 278056 443550 278438 443578
rect 278792 443550 279266 443578
rect 279620 443550 280002 443578
rect 280356 443550 280830 443578
rect 281566 443550 281764 443578
rect 281920 443578 281948 447034
rect 283024 443578 283052 454718
rect 284312 447098 284340 476342
rect 285680 476332 285732 476338
rect 285680 476274 285732 476280
rect 284392 474088 284444 474094
rect 284392 474030 284444 474036
rect 283564 447092 283616 447098
rect 283564 447034 283616 447040
rect 284300 447092 284352 447098
rect 284300 447034 284352 447040
rect 283576 443578 283604 447034
rect 284404 443578 284432 474030
rect 285692 447098 285720 476274
rect 288440 476264 288492 476270
rect 285770 476232 285826 476241
rect 285770 476167 285826 476176
rect 287058 476232 287114 476241
rect 288440 476206 288492 476212
rect 289910 476232 289966 476241
rect 287058 476167 287114 476176
rect 285784 463010 285812 476167
rect 285772 463004 285824 463010
rect 285772 462946 285824 462952
rect 285772 461712 285824 461718
rect 285772 461654 285824 461660
rect 285784 460934 285812 461654
rect 285784 460906 285904 460934
rect 285036 447092 285088 447098
rect 285036 447034 285088 447040
rect 285680 447092 285732 447098
rect 285680 447034 285732 447040
rect 285048 443578 285076 447034
rect 285876 443578 285904 460906
rect 287072 457570 287100 476167
rect 287060 457564 287112 457570
rect 287060 457506 287112 457512
rect 287336 453416 287388 453422
rect 287336 453358 287388 453364
rect 286692 447092 286744 447098
rect 286692 447034 286744 447040
rect 286704 443578 286732 447034
rect 287348 443578 287376 453358
rect 288452 443578 288480 476206
rect 289820 476196 289872 476202
rect 289910 476167 289966 476176
rect 289820 476138 289872 476144
rect 288808 451920 288860 451926
rect 288808 451862 288860 451868
rect 288820 443578 288848 451862
rect 289832 443578 289860 476138
rect 289924 458930 289952 476167
rect 289912 458924 289964 458930
rect 289912 458866 289964 458872
rect 290464 454708 290516 454714
rect 290464 454650 290516 454656
rect 290476 443578 290504 454650
rect 291212 443578 291240 476682
rect 292578 476232 292634 476241
rect 292578 476167 292634 476176
rect 295430 476232 295486 476241
rect 295430 476167 295486 476176
rect 298190 476232 298246 476241
rect 298190 476167 298246 476176
rect 300950 476232 301006 476241
rect 300950 476167 301006 476176
rect 292592 453354 292620 476167
rect 295340 467220 295392 467226
rect 295340 467162 295392 467168
rect 292580 453348 292632 453354
rect 292580 453290 292632 453296
rect 294328 451920 294380 451926
rect 294328 451862 294380 451868
rect 293132 446276 293184 446282
rect 293132 446218 293184 446224
rect 292396 446208 292448 446214
rect 292396 446150 292448 446156
rect 281920 443550 282302 443578
rect 283024 443550 283130 443578
rect 283576 443550 283866 443578
rect 284404 443550 284694 443578
rect 285048 443550 285430 443578
rect 285876 443550 286258 443578
rect 286704 443550 286994 443578
rect 287348 443550 287730 443578
rect 288452 443550 288558 443578
rect 288820 443550 289294 443578
rect 289832 443550 290122 443578
rect 290476 443550 290858 443578
rect 291212 443550 291686 443578
rect 292408 443564 292436 446150
rect 293144 443564 293172 446218
rect 293960 445868 294012 445874
rect 293960 445810 294012 445816
rect 293972 443564 294000 445810
rect 294340 443578 294368 451862
rect 295352 451274 295380 467162
rect 295444 460290 295472 476167
rect 298100 474088 298152 474094
rect 298100 474030 298152 474036
rect 295432 460284 295484 460290
rect 295432 460226 295484 460232
rect 296720 453348 296772 453354
rect 296720 453290 296772 453296
rect 295352 451246 295840 451274
rect 295524 444780 295576 444786
rect 295524 444722 295576 444728
rect 294340 443550 294722 443578
rect 295536 443564 295564 444722
rect 295812 443578 295840 451246
rect 296732 443578 296760 453290
rect 298112 443578 298140 474030
rect 298204 464438 298232 476167
rect 300860 469940 300912 469946
rect 300860 469882 300912 469888
rect 298192 464432 298244 464438
rect 298192 464374 298244 464380
rect 298928 454708 298980 454714
rect 298928 454650 298980 454656
rect 298940 443578 298968 454650
rect 300124 444848 300176 444854
rect 300124 444790 300176 444796
rect 295812 443550 296286 443578
rect 296732 443550 297114 443578
rect 298112 443550 298678 443578
rect 298940 443550 299414 443578
rect 300136 443564 300164 444790
rect 300872 443578 300900 469882
rect 300964 465798 300992 476167
rect 302252 476134 302280 476847
rect 305012 476678 305040 476983
rect 305000 476672 305052 476678
rect 305000 476614 305052 476620
rect 307772 476610 307800 476983
rect 307760 476604 307812 476610
rect 307760 476546 307812 476552
rect 302240 476128 302292 476134
rect 302240 476070 302292 476076
rect 300952 465792 301004 465798
rect 300952 465734 301004 465740
rect 307760 464432 307812 464438
rect 307760 464374 307812 464380
rect 307772 460934 307800 464374
rect 309152 460934 309180 478246
rect 314752 478236 314804 478242
rect 314752 478178 314804 478184
rect 310518 476912 310574 476921
rect 310518 476847 310574 476856
rect 310532 476542 310560 476847
rect 310520 476536 310572 476542
rect 310520 476478 310572 476484
rect 313278 476504 313334 476513
rect 313278 476439 313280 476448
rect 313332 476439 313334 476448
rect 314658 476504 314714 476513
rect 314658 476439 314714 476448
rect 313280 476410 313332 476416
rect 314672 476406 314700 476439
rect 314660 476400 314712 476406
rect 314660 476342 314712 476348
rect 314764 470594 314792 478178
rect 346492 478168 346544 478174
rect 346492 478110 346544 478116
rect 322938 476912 322994 476921
rect 322938 476847 322994 476856
rect 325790 476912 325846 476921
rect 325790 476847 325846 476856
rect 317418 476368 317474 476377
rect 317418 476303 317420 476312
rect 317472 476303 317474 476312
rect 320178 476368 320234 476377
rect 320178 476303 320234 476312
rect 317420 476274 317472 476280
rect 320192 476270 320220 476303
rect 320180 476264 320232 476270
rect 320180 476206 320232 476212
rect 322952 476202 322980 476847
rect 325804 476746 325832 476847
rect 325792 476740 325844 476746
rect 325792 476682 325844 476688
rect 322940 476196 322992 476202
rect 322940 476138 322992 476144
rect 331220 474768 331272 474774
rect 331220 474710 331272 474716
rect 324320 474020 324372 474026
rect 324320 473962 324372 473968
rect 314672 470566 314792 470594
rect 307772 460906 308352 460934
rect 309152 460906 309824 460934
rect 306380 458924 306432 458930
rect 306380 458866 306432 458872
rect 303712 457564 303764 457570
rect 303712 457506 303764 457512
rect 301320 456136 301372 456142
rect 301320 456078 301372 456084
rect 301332 443578 301360 456078
rect 303252 449336 303304 449342
rect 303252 449278 303304 449284
rect 302516 445800 302568 445806
rect 302516 445742 302568 445748
rect 300872 443550 300978 443578
rect 301332 443550 301714 443578
rect 302528 443564 302556 445742
rect 303264 443564 303292 449278
rect 303724 443578 303752 457506
rect 305552 449472 305604 449478
rect 305552 449414 305604 449420
rect 304816 446344 304868 446350
rect 304816 446286 304868 446292
rect 303724 443550 304106 443578
rect 304828 443564 304856 446286
rect 305564 443564 305592 449414
rect 306392 443564 306420 458866
rect 307944 449608 307996 449614
rect 307944 449550 307996 449556
rect 307116 446480 307168 446486
rect 307116 446422 307168 446428
rect 307128 443564 307156 446422
rect 307956 443564 307984 449550
rect 308324 443578 308352 460906
rect 309508 443760 309560 443766
rect 309508 443702 309560 443708
rect 308324 443550 308706 443578
rect 309520 443564 309548 443702
rect 309796 443578 309824 460906
rect 313372 446684 313424 446690
rect 313372 446626 313424 446632
rect 312544 446616 312596 446622
rect 312544 446558 312596 446564
rect 310980 446548 311032 446554
rect 310980 446490 311032 446496
rect 309796 443550 310270 443578
rect 310992 443564 311020 446490
rect 311808 446412 311860 446418
rect 311808 446354 311860 446360
rect 311164 445800 311216 445806
rect 311164 445742 311216 445748
rect 311176 445058 311204 445742
rect 311164 445052 311216 445058
rect 311164 444994 311216 445000
rect 311820 443564 311848 446354
rect 312556 443564 312584 446558
rect 313384 443564 313412 446626
rect 314384 443692 314436 443698
rect 314384 443634 314436 443640
rect 314396 443578 314424 443634
rect 314134 443550 314424 443578
rect 314672 443578 314700 470566
rect 317420 468512 317472 468518
rect 317420 468454 317472 468460
rect 320180 468512 320232 468518
rect 320180 468454 320232 468460
rect 314752 465724 314804 465730
rect 314752 465666 314804 465672
rect 314764 460934 314792 465666
rect 317432 460934 317460 468454
rect 318800 465724 318852 465730
rect 318800 465666 318852 465672
rect 314764 460906 315344 460934
rect 317432 460906 317552 460934
rect 315316 443578 315344 460906
rect 317236 449540 317288 449546
rect 317236 449482 317288 449488
rect 316408 445800 316460 445806
rect 316408 445742 316460 445748
rect 314672 443550 314962 443578
rect 315316 443550 315698 443578
rect 316420 443564 316448 445742
rect 317248 443564 317276 449482
rect 317524 443578 317552 460906
rect 317524 443550 317998 443578
rect 318812 443564 318840 465666
rect 320192 460934 320220 468454
rect 321560 467152 321612 467158
rect 321560 467094 321612 467100
rect 321572 460934 321600 467094
rect 324332 460934 324360 473962
rect 328460 472660 328512 472666
rect 328460 472602 328512 472608
rect 327080 469872 327132 469878
rect 327080 469814 327132 469820
rect 325700 461644 325752 461650
rect 325700 461586 325752 461592
rect 320192 460906 320680 460934
rect 321572 460906 322336 460934
rect 324332 460906 324544 460934
rect 319536 449404 319588 449410
rect 319536 449346 319588 449352
rect 319548 443564 319576 449346
rect 320364 447908 320416 447914
rect 320364 447850 320416 447856
rect 320376 443564 320404 447850
rect 320652 443578 320680 460906
rect 321836 449268 321888 449274
rect 321836 449210 321888 449216
rect 320652 443550 321126 443578
rect 321848 443564 321876 449210
rect 322308 443578 322336 460906
rect 322940 460284 322992 460290
rect 322940 460226 322992 460232
rect 322952 443578 322980 460226
rect 323768 456068 323820 456074
rect 323768 456010 323820 456016
rect 323780 443578 323808 456010
rect 324516 443578 324544 460906
rect 325712 443578 325740 461586
rect 326528 449200 326580 449206
rect 326528 449142 326580 449148
rect 322308 443550 322690 443578
rect 322952 443550 323426 443578
rect 323780 443550 324254 443578
rect 324516 443550 324990 443578
rect 325712 443550 325818 443578
rect 326540 443564 326568 449142
rect 327092 443578 327120 469814
rect 328472 460934 328500 472602
rect 331232 460934 331260 474710
rect 332600 462392 332652 462398
rect 332600 462334 332652 462340
rect 332612 460934 332640 462334
rect 328472 460906 329328 460934
rect 331232 460906 331536 460934
rect 332612 460906 333192 460934
rect 328092 450696 328144 450702
rect 328092 450638 328144 450644
rect 327092 443550 327290 443578
rect 328104 443564 328132 450638
rect 328828 450628 328880 450634
rect 328828 450570 328880 450576
rect 328840 443564 328868 450570
rect 329300 443578 329328 460906
rect 331220 450560 331272 450566
rect 331220 450502 331272 450508
rect 330392 447908 330444 447914
rect 330392 447850 330444 447856
rect 329300 443550 329682 443578
rect 330404 443564 330432 447850
rect 331232 443564 331260 450502
rect 331508 443578 331536 460906
rect 332784 448112 332836 448118
rect 332784 448054 332836 448060
rect 331508 443550 331982 443578
rect 332796 443564 332824 448054
rect 333164 443578 333192 460906
rect 335084 448180 335136 448186
rect 335084 448122 335136 448128
rect 333980 445800 334032 445806
rect 333980 445742 334032 445748
rect 333992 445126 334020 445742
rect 333980 445120 334032 445126
rect 333980 445062 334032 445068
rect 334256 444440 334308 444446
rect 334256 444382 334308 444388
rect 333164 443550 333546 443578
rect 334268 443564 334296 444382
rect 335096 443564 335124 448122
rect 342076 448044 342128 448050
rect 342076 447986 342128 447992
rect 339684 446752 339736 446758
rect 339684 446694 339736 446700
rect 337384 446684 337436 446690
rect 337384 446626 337436 446632
rect 336648 445256 336700 445262
rect 336648 445198 336700 445204
rect 335556 443562 335846 443578
rect 336660 443564 336688 445198
rect 337396 443564 337424 446626
rect 338212 446072 338264 446078
rect 338212 446014 338264 446020
rect 338224 443564 338252 446014
rect 338948 445188 339000 445194
rect 338948 445130 339000 445136
rect 338960 443564 338988 445130
rect 339696 443564 339724 446694
rect 341248 444984 341300 444990
rect 341248 444926 341300 444932
rect 341260 443564 341288 444926
rect 342088 443564 342116 447986
rect 344376 447976 344428 447982
rect 344376 447918 344428 447924
rect 343640 444712 343692 444718
rect 343640 444654 343692 444660
rect 343652 443564 343680 444654
rect 344388 443564 344416 447918
rect 345112 446140 345164 446146
rect 345112 446082 345164 446088
rect 345124 443564 345152 446082
rect 345940 444644 345992 444650
rect 345940 444586 345992 444592
rect 345952 443564 345980 444586
rect 346504 443578 346532 478110
rect 347872 471300 347924 471306
rect 347872 471242 347924 471248
rect 347884 460934 347912 471242
rect 350540 464364 350592 464370
rect 350540 464306 350592 464312
rect 347884 460906 348648 460934
rect 347504 446004 347556 446010
rect 347504 445946 347556 445952
rect 335544 443556 335846 443562
rect 335596 443550 335846 443556
rect 346504 443550 346702 443578
rect 347516 443564 347544 445946
rect 348240 444576 348292 444582
rect 348240 444518 348292 444524
rect 348252 443564 348280 444518
rect 348620 443578 348648 460906
rect 350552 447098 350580 464306
rect 350632 460216 350684 460222
rect 350632 460158 350684 460164
rect 350540 447092 350592 447098
rect 350540 447034 350592 447040
rect 349804 446820 349856 446826
rect 349804 446762 349856 446768
rect 348620 443550 349094 443578
rect 349816 443564 349844 446762
rect 350644 443578 350672 460158
rect 351920 458856 351972 458862
rect 351920 458798 351972 458804
rect 351092 447092 351144 447098
rect 351092 447034 351144 447040
rect 350566 443550 350672 443578
rect 351104 443578 351132 447034
rect 351932 443578 351960 458798
rect 352472 457496 352524 457502
rect 352472 457438 352524 457444
rect 352484 443578 352512 457438
rect 353668 447840 353720 447846
rect 353668 447782 353720 447788
rect 351104 443550 351394 443578
rect 351932 443550 352130 443578
rect 352484 443550 352958 443578
rect 353680 443564 353708 447782
rect 357452 446758 357480 700266
rect 357440 446752 357492 446758
rect 357440 446694 357492 446700
rect 357544 446554 357572 700402
rect 357636 478310 357664 700538
rect 358912 700528 358964 700534
rect 358912 700470 358964 700476
rect 358820 700392 358872 700398
rect 358820 700334 358872 700340
rect 357624 478304 357676 478310
rect 357624 478246 357676 478252
rect 358832 446622 358860 700334
rect 358924 446690 358952 700470
rect 360844 670744 360896 670750
rect 360844 670686 360896 670692
rect 359464 563100 359516 563106
rect 359464 563042 359516 563048
rect 359476 451926 359504 563042
rect 360856 454714 360884 670686
rect 363604 590708 363656 590714
rect 363604 590650 363656 590656
rect 363616 460290 363644 590650
rect 364352 464438 364380 702406
rect 371884 700324 371936 700330
rect 371884 700266 371936 700272
rect 369124 696992 369176 696998
rect 369124 696934 369176 696940
rect 367744 576904 367796 576910
rect 367744 576846 367796 576852
rect 367756 467226 367784 576846
rect 367744 467220 367796 467226
rect 367744 467162 367796 467168
rect 364340 464432 364392 464438
rect 364340 464374 364392 464380
rect 363604 460284 363656 460290
rect 363604 460226 363656 460232
rect 360844 454708 360896 454714
rect 360844 454650 360896 454656
rect 359464 451920 359516 451926
rect 359464 451862 359516 451868
rect 369136 450702 369164 696934
rect 371896 456142 371924 700266
rect 373264 643136 373316 643142
rect 373264 643078 373316 643084
rect 373276 461650 373304 643078
rect 377404 630692 377456 630698
rect 377404 630634 377456 630640
rect 377416 474094 377444 630634
rect 378784 616888 378836 616894
rect 378784 616830 378836 616836
rect 377404 474088 377456 474094
rect 377404 474030 377456 474036
rect 373264 461644 373316 461650
rect 373264 461586 373316 461592
rect 371884 456136 371936 456142
rect 371884 456078 371936 456084
rect 378796 453354 378824 616830
rect 378784 453348 378836 453354
rect 378784 453290 378836 453296
rect 369124 450696 369176 450702
rect 369124 450638 369176 450644
rect 397472 448186 397500 703520
rect 412652 449614 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 699718 429884 703520
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 428476 458930 428504 699654
rect 428464 458924 428516 458930
rect 428464 458866 428516 458872
rect 412640 449608 412692 449614
rect 412640 449550 412692 449556
rect 397460 448180 397512 448186
rect 397460 448122 397512 448128
rect 462332 448118 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 449478 477540 702406
rect 482284 484424 482336 484430
rect 482284 484366 482336 484372
rect 482296 465730 482324 484366
rect 482284 465724 482336 465730
rect 482284 465666 482336 465672
rect 494072 457570 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 500224 536852 500276 536858
rect 500224 536794 500276 536800
rect 500236 468518 500264 536794
rect 500224 468512 500276 468518
rect 500224 468454 500276 468460
rect 494060 457564 494112 457570
rect 494060 457506 494112 457512
rect 477500 449472 477552 449478
rect 477500 449414 477552 449420
rect 462320 448112 462372 448118
rect 462320 448054 462372 448060
rect 527192 447914 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 449342 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580276 469946 580304 683839
rect 580264 469940 580316 469946
rect 580264 469882 580316 469888
rect 542360 449336 542412 449342
rect 542360 449278 542412 449284
rect 527180 447908 527232 447914
rect 527180 447850 527232 447856
rect 358912 446684 358964 446690
rect 358912 446626 358964 446632
rect 358820 446616 358872 446622
rect 358820 446558 358872 446564
rect 357532 446548 357584 446554
rect 357532 446490 357584 446496
rect 364984 446480 365036 446486
rect 364984 446422 365036 446428
rect 362224 446412 362276 446418
rect 362224 446354 362276 446360
rect 359924 445936 359976 445942
rect 359924 445878 359976 445884
rect 355968 444916 356020 444922
rect 355968 444858 356020 444864
rect 355980 443564 356008 444858
rect 358360 444508 358412 444514
rect 358360 444450 358412 444456
rect 358372 443564 358400 444450
rect 359936 443564 359964 445878
rect 335544 443498 335596 443504
rect 340236 443488 340288 443494
rect 340288 443436 340538 443442
rect 340236 443430 340538 443436
rect 340248 443414 340538 443430
rect 342456 443426 342838 443442
rect 342444 443420 342838 443426
rect 342496 443414 342838 443420
rect 342444 443362 342496 443368
rect 354220 443352 354272 443358
rect 354272 443300 354522 443306
rect 354220 443294 354522 443300
rect 354232 443278 354522 443294
rect 354968 443290 355258 443306
rect 354956 443284 355258 443290
rect 355008 443278 355258 443284
rect 354956 443226 355008 443232
rect 298008 443216 298060 443222
rect 297850 443164 298008 443170
rect 297850 443158 298060 443164
rect 297850 443142 298048 443158
rect 356440 443154 356822 443170
rect 356428 443148 356822 443154
rect 356480 443142 356822 443148
rect 356428 443090 356480 443096
rect 357440 443080 357492 443086
rect 358820 443080 358872 443086
rect 357492 443028 357558 443034
rect 357440 443022 357558 443028
rect 358872 443028 359122 443034
rect 358820 443022 359122 443028
rect 357452 443006 357558 443022
rect 358832 443006 359122 443022
rect 360686 443006 361160 443034
rect 229836 442264 229888 442270
rect 229836 442206 229888 442212
rect 229744 410576 229796 410582
rect 229744 410518 229796 410524
rect 228640 398812 228692 398818
rect 228640 398754 228692 398760
rect 228548 372564 228600 372570
rect 228548 372506 228600 372512
rect 261220 310554 261418 310570
rect 261024 310548 261076 310554
rect 261024 310490 261076 310496
rect 261208 310548 261418 310554
rect 261260 310542 261418 310548
rect 266386 310554 266584 310570
rect 291672 310554 291870 310570
rect 292960 310554 293158 310570
rect 301240 310554 301438 310570
rect 310808 310554 311006 310570
rect 327552 310554 327750 310570
rect 266386 310548 266596 310554
rect 266386 310542 266544 310548
rect 261208 310490 261260 310496
rect 266544 310490 266596 310496
rect 266728 310548 266780 310554
rect 266728 310490 266780 310496
rect 291476 310548 291528 310554
rect 291476 310490 291528 310496
rect 291660 310548 291870 310554
rect 291712 310542 291870 310548
rect 292764 310548 292816 310554
rect 291660 310490 291712 310496
rect 292764 310490 292816 310496
rect 292948 310548 293158 310554
rect 293000 310542 293158 310548
rect 300860 310548 300912 310554
rect 292948 310490 293000 310496
rect 300860 310490 300912 310496
rect 301228 310548 301438 310554
rect 301280 310542 301438 310548
rect 310612 310548 310664 310554
rect 301228 310490 301280 310496
rect 310612 310490 310664 310496
rect 310796 310548 311006 310554
rect 310848 310542 311006 310548
rect 327356 310548 327408 310554
rect 310796 310490 310848 310496
rect 327356 310490 327408 310496
rect 327540 310548 327750 310554
rect 327592 310542 327750 310548
rect 353326 310554 353524 310570
rect 353326 310548 353536 310554
rect 353326 310542 353484 310548
rect 327540 310490 327592 310496
rect 353484 310490 353536 310496
rect 353668 310548 353720 310554
rect 356178 310542 356376 310570
rect 353668 310490 353720 310496
rect 229652 309120 229704 309126
rect 229652 309062 229704 309068
rect 229664 308718 229692 309062
rect 229744 308984 229796 308990
rect 229744 308926 229796 308932
rect 229652 308712 229704 308718
rect 229652 308654 229704 308660
rect 229756 308650 229784 308926
rect 229744 308644 229796 308650
rect 229744 308586 229796 308592
rect 229744 307828 229796 307834
rect 229744 307770 229796 307776
rect 229192 306332 229244 306338
rect 229192 306274 229244 306280
rect 228456 293956 228508 293962
rect 228456 293898 228508 293904
rect 229204 247722 229232 306274
rect 229756 262886 229784 307770
rect 230124 307086 230152 310420
rect 230112 307080 230164 307086
rect 230112 307022 230164 307028
rect 230308 306338 230336 310420
rect 230296 306332 230348 306338
rect 230296 306274 230348 306280
rect 230492 304298 230520 310420
rect 230768 306354 230796 310420
rect 230952 307834 230980 310420
rect 230940 307828 230992 307834
rect 230940 307770 230992 307776
rect 230768 306326 231072 306354
rect 230940 306264 230992 306270
rect 230940 306206 230992 306212
rect 230848 305992 230900 305998
rect 230848 305934 230900 305940
rect 230480 304292 230532 304298
rect 230480 304234 230532 304240
rect 230664 304156 230716 304162
rect 230664 304098 230716 304104
rect 230676 287706 230704 304098
rect 230664 287700 230716 287706
rect 230664 287642 230716 287648
rect 229744 262880 229796 262886
rect 229744 262822 229796 262828
rect 229192 247716 229244 247722
rect 229192 247658 229244 247664
rect 228364 246356 228416 246362
rect 228364 246298 228416 246304
rect 230860 244934 230888 305934
rect 230952 274038 230980 306206
rect 231044 300150 231072 306326
rect 231136 305998 231164 310420
rect 231124 305992 231176 305998
rect 231124 305934 231176 305940
rect 231412 302938 231440 310420
rect 231596 306270 231624 310420
rect 231584 306264 231636 306270
rect 231584 306206 231636 306212
rect 231780 304162 231808 310420
rect 232056 308582 232084 310420
rect 232044 308576 232096 308582
rect 232044 308518 232096 308524
rect 232044 306400 232096 306406
rect 232044 306342 232096 306348
rect 231952 306332 232004 306338
rect 231952 306274 232004 306280
rect 231768 304156 231820 304162
rect 231768 304098 231820 304104
rect 231400 302932 231452 302938
rect 231400 302874 231452 302880
rect 231032 300144 231084 300150
rect 231032 300086 231084 300092
rect 230940 274032 230992 274038
rect 230940 273974 230992 273980
rect 231964 258738 231992 306274
rect 232056 283626 232084 306342
rect 232240 302234 232268 310420
rect 232148 302206 232268 302234
rect 232148 289134 232176 302206
rect 232424 296714 232452 310420
rect 232516 310406 232714 310434
rect 232516 306338 232544 310406
rect 232884 308786 232912 310420
rect 232976 310406 233174 310434
rect 232872 308780 232924 308786
rect 232872 308722 232924 308728
rect 232976 306406 233004 310406
rect 232964 306400 233016 306406
rect 232964 306342 233016 306348
rect 232504 306332 232556 306338
rect 232504 306274 232556 306280
rect 232240 296686 232452 296714
rect 232136 289128 232188 289134
rect 232136 289070 232188 289076
rect 232044 283620 232096 283626
rect 232044 283562 232096 283568
rect 231952 258732 232004 258738
rect 231952 258674 232004 258680
rect 232240 249082 232268 296686
rect 233344 251870 233372 310420
rect 233528 306746 233556 310420
rect 233620 310406 233818 310434
rect 233516 306740 233568 306746
rect 233516 306682 233568 306688
rect 233516 306536 233568 306542
rect 233516 306478 233568 306484
rect 233424 304292 233476 304298
rect 233424 304234 233476 304240
rect 233436 261526 233464 304234
rect 233528 275330 233556 306478
rect 233620 304298 233648 310406
rect 233608 304292 233660 304298
rect 233608 304234 233660 304240
rect 233988 302234 234016 310420
rect 233620 302206 234016 302234
rect 233620 282198 233648 302206
rect 234172 296714 234200 310420
rect 234448 308446 234476 310420
rect 234632 308854 234660 310420
rect 234620 308848 234672 308854
rect 234620 308790 234672 308796
rect 234436 308440 234488 308446
rect 234436 308382 234488 308388
rect 234712 306468 234764 306474
rect 234712 306410 234764 306416
rect 233712 296686 234200 296714
rect 233608 282192 233660 282198
rect 233608 282134 233660 282140
rect 233516 275324 233568 275330
rect 233516 275266 233568 275272
rect 233424 261520 233476 261526
rect 233424 261462 233476 261468
rect 233332 251864 233384 251870
rect 233332 251806 233384 251812
rect 233712 250510 233740 296686
rect 234724 279478 234752 306410
rect 234816 280838 234844 310420
rect 234908 310406 235106 310434
rect 234908 294642 234936 310406
rect 235276 308514 235304 310420
rect 235368 310406 235566 310434
rect 235264 308508 235316 308514
rect 235264 308450 235316 308456
rect 235368 306474 235396 310406
rect 235356 306468 235408 306474
rect 235356 306410 235408 306416
rect 235736 306354 235764 310420
rect 235920 308990 235948 310420
rect 236104 310406 236210 310434
rect 235908 308984 235960 308990
rect 235908 308926 235960 308932
rect 235816 308780 235868 308786
rect 235816 308722 235868 308728
rect 235000 306326 235764 306354
rect 234896 294636 234948 294642
rect 234896 294578 234948 294584
rect 234804 280832 234856 280838
rect 234804 280774 234856 280780
rect 234712 279472 234764 279478
rect 234712 279414 234764 279420
rect 235000 253230 235028 306326
rect 235828 302234 235856 308722
rect 235276 302206 235856 302234
rect 235276 282266 235304 302206
rect 235264 282260 235316 282266
rect 235264 282202 235316 282208
rect 236104 278050 236132 310406
rect 236380 306354 236408 310420
rect 236564 309126 236592 310420
rect 236656 310406 236854 310434
rect 236552 309120 236604 309126
rect 236552 309062 236604 309068
rect 236184 306332 236236 306338
rect 236184 306274 236236 306280
rect 236288 306326 236408 306354
rect 236196 284986 236224 306274
rect 236288 291854 236316 306326
rect 236656 306082 236684 310406
rect 236828 308508 236880 308514
rect 236828 308450 236880 308456
rect 236736 307828 236788 307834
rect 236736 307770 236788 307776
rect 236380 306054 236684 306082
rect 236276 291848 236328 291854
rect 236276 291790 236328 291796
rect 236184 284980 236236 284986
rect 236184 284922 236236 284928
rect 236092 278044 236144 278050
rect 236092 277986 236144 277992
rect 236380 276690 236408 306054
rect 236644 305380 236696 305386
rect 236644 305322 236696 305328
rect 236368 276684 236420 276690
rect 236368 276626 236420 276632
rect 236656 254590 236684 305322
rect 236748 275398 236776 307770
rect 236840 305386 236868 308450
rect 237024 306338 237052 310420
rect 237208 309058 237236 310420
rect 237484 309134 237512 310420
rect 237668 309134 237696 310420
rect 237392 309106 237512 309134
rect 237576 309106 237696 309134
rect 237196 309052 237248 309058
rect 237196 308994 237248 309000
rect 237012 306332 237064 306338
rect 237012 306274 237064 306280
rect 236828 305380 236880 305386
rect 236828 305322 236880 305328
rect 237392 301510 237420 309106
rect 237472 306264 237524 306270
rect 237472 306206 237524 306212
rect 237576 306218 237604 309106
rect 237944 306270 237972 310420
rect 238024 308440 238076 308446
rect 238024 308382 238076 308388
rect 238036 307170 238064 308382
rect 238128 307834 238156 310420
rect 238206 308408 238262 308417
rect 238206 308343 238262 308352
rect 238116 307828 238168 307834
rect 238116 307770 238168 307776
rect 238036 307142 238156 307170
rect 238024 307080 238076 307086
rect 238024 307022 238076 307028
rect 237932 306264 237984 306270
rect 237380 301504 237432 301510
rect 237380 301446 237432 301452
rect 236736 275392 236788 275398
rect 236736 275334 236788 275340
rect 237484 260166 237512 306206
rect 237576 306190 237696 306218
rect 237932 306206 237984 306212
rect 237564 306128 237616 306134
rect 237564 306070 237616 306076
rect 237576 286346 237604 306070
rect 237668 290494 237696 306190
rect 237748 306196 237800 306202
rect 237748 306138 237800 306144
rect 237656 290488 237708 290494
rect 237656 290430 237708 290436
rect 237564 286340 237616 286346
rect 237564 286282 237616 286288
rect 237472 260160 237524 260166
rect 237472 260102 237524 260108
rect 236644 254584 236696 254590
rect 236644 254526 236696 254532
rect 234988 253224 235040 253230
rect 234988 253166 235040 253172
rect 233700 250504 233752 250510
rect 233700 250446 233752 250452
rect 232228 249076 232280 249082
rect 232228 249018 232280 249024
rect 230848 244928 230900 244934
rect 230848 244870 230900 244876
rect 236736 170400 236788 170406
rect 236736 170342 236788 170348
rect 99286 168056 99342 168065
rect 99286 167991 99342 168000
rect 153658 159896 153714 159905
rect 153658 159831 153714 159840
rect 156050 159896 156106 159905
rect 156050 159831 156106 159840
rect 160926 159896 160982 159905
rect 160926 159831 160982 159840
rect 175922 159896 175978 159905
rect 175922 159831 175978 159840
rect 153672 158914 153700 159831
rect 156064 158982 156092 159831
rect 160940 159050 160968 159831
rect 165986 159624 166042 159633
rect 165986 159559 166042 159568
rect 166000 159118 166028 159559
rect 165988 159112 166040 159118
rect 165988 159054 166040 159060
rect 160928 159044 160980 159050
rect 160928 158986 160980 158992
rect 156052 158976 156104 158982
rect 156052 158918 156104 158924
rect 153660 158908 153712 158914
rect 153660 158850 153712 158856
rect 168288 158840 168340 158846
rect 168288 158782 168340 158788
rect 128728 158704 128780 158710
rect 116214 158672 116270 158681
rect 116214 158607 116270 158616
rect 118238 158672 118294 158681
rect 118238 158607 118294 158616
rect 119894 158672 119950 158681
rect 119894 158607 119950 158616
rect 120630 158672 120686 158681
rect 120630 158607 120686 158616
rect 121918 158672 121974 158681
rect 121918 158607 121974 158616
rect 126518 158672 126574 158681
rect 126518 158607 126520 158616
rect 116228 157350 116256 158607
rect 117226 158128 117282 158137
rect 117282 158086 117360 158114
rect 117226 158063 117282 158072
rect 116216 157344 116268 157350
rect 116216 157286 116268 157292
rect 117332 156194 117360 158086
rect 118252 157282 118280 158607
rect 119908 157758 119936 158607
rect 120644 158506 120672 158607
rect 121932 158574 121960 158607
rect 126572 158607 126574 158616
rect 127622 158672 127678 158681
rect 127622 158607 127678 158616
rect 128726 158672 128728 158681
rect 168300 158681 168328 158782
rect 175936 158778 175964 159831
rect 236748 159662 236776 170342
rect 236736 159656 236788 159662
rect 236736 159598 236788 159604
rect 234620 159452 234672 159458
rect 234620 159394 234672 159400
rect 220820 159384 220872 159390
rect 200118 159352 200174 159361
rect 220820 159326 220872 159332
rect 200118 159287 200174 159296
rect 175924 158772 175976 158778
rect 175924 158714 175976 158720
rect 128780 158672 128782 158681
rect 128726 158607 128782 158616
rect 130566 158672 130622 158681
rect 130566 158607 130622 158616
rect 131302 158672 131358 158681
rect 131302 158607 131358 158616
rect 132406 158672 132462 158681
rect 132406 158607 132462 158616
rect 133510 158672 133566 158681
rect 133510 158607 133566 158616
rect 139306 158672 139362 158681
rect 139306 158607 139362 158616
rect 159638 158672 159694 158681
rect 159638 158607 159694 158616
rect 168286 158672 168342 158681
rect 168286 158607 168342 158616
rect 188710 158672 188766 158681
rect 188710 158607 188766 158616
rect 126520 158578 126572 158584
rect 121920 158568 121972 158574
rect 121920 158510 121972 158516
rect 120632 158500 120684 158506
rect 120632 158442 120684 158448
rect 127636 158370 127664 158607
rect 127624 158364 127676 158370
rect 127624 158306 127676 158312
rect 123942 158264 123998 158273
rect 123942 158199 123998 158208
rect 119896 157752 119948 157758
rect 119896 157694 119948 157700
rect 118240 157276 118292 157282
rect 118240 157218 118292 157224
rect 123956 156330 123984 158199
rect 130580 157622 130608 158607
rect 131316 158234 131344 158607
rect 132420 158302 132448 158607
rect 132408 158296 132460 158302
rect 132408 158238 132460 158244
rect 131304 158228 131356 158234
rect 131304 158170 131356 158176
rect 133524 158098 133552 158607
rect 135902 158536 135958 158545
rect 135902 158471 135958 158480
rect 137006 158536 137062 158545
rect 137006 158471 137062 158480
rect 138386 158536 138442 158545
rect 138386 158471 138442 158480
rect 134614 158264 134670 158273
rect 134614 158199 134670 158208
rect 133512 158092 133564 158098
rect 133512 158034 133564 158040
rect 130568 157616 130620 157622
rect 124770 157584 124826 157593
rect 130568 157558 130620 157564
rect 124770 157519 124826 157528
rect 123944 156324 123996 156330
rect 123944 156266 123996 156272
rect 117320 156188 117372 156194
rect 117320 156130 117372 156136
rect 124784 154902 124812 157519
rect 125414 157448 125470 157457
rect 125414 157383 125470 157392
rect 133694 157448 133750 157457
rect 133694 157383 133750 157392
rect 124772 154896 124824 154902
rect 124772 154838 124824 154844
rect 125428 154562 125456 157383
rect 125600 156664 125652 156670
rect 125600 156606 125652 156612
rect 125416 154556 125468 154562
rect 125416 154498 125468 154504
rect 121460 141432 121512 141438
rect 121460 141374 121512 141380
rect 114560 140072 114612 140078
rect 114560 140014 114612 140020
rect 107660 137284 107712 137290
rect 107660 137226 107712 137232
rect 103520 135924 103572 135930
rect 103520 135866 103572 135872
rect 100760 130416 100812 130422
rect 100760 130358 100812 130364
rect 99380 90364 99432 90370
rect 99380 90306 99432 90312
rect 99392 16574 99420 90306
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 97264 3664 97316 3670
rect 97264 3606 97316 3612
rect 97184 3454 97488 3482
rect 97460 480 97488 3454
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 130358
rect 102140 22772 102192 22778
rect 102140 22714 102192 22720
rect 102152 3398 102180 22714
rect 103532 16574 103560 135866
rect 106280 91792 106332 91798
rect 106280 91734 106332 91740
rect 106292 16574 106320 91734
rect 107672 16574 107700 137226
rect 110420 131776 110472 131782
rect 110420 131718 110472 131724
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102232 3664 102284 3670
rect 102232 3606 102284 3612
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 3606
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 11756 105780 11762
rect 105728 11698 105780 11704
rect 105740 480 105768 11698
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109316 8968 109368 8974
rect 109316 8910 109368 8916
rect 109328 480 109356 8910
rect 110432 3398 110460 131718
rect 111800 94512 111852 94518
rect 111800 94454 111852 94460
rect 110512 24132 110564 24138
rect 110512 24074 110564 24080
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 24074
rect 111812 16574 111840 94454
rect 113180 86284 113232 86290
rect 113180 86226 113232 86232
rect 113192 16574 113220 86226
rect 114572 16574 114600 140014
rect 118700 102808 118752 102814
rect 118700 102750 118752 102756
rect 115940 93152 115992 93158
rect 115940 93094 115992 93100
rect 115952 16574 115980 93094
rect 117320 87644 117372 87650
rect 117320 87586 117372 87592
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 87586
rect 118712 16574 118740 102750
rect 121472 16574 121500 141374
rect 118712 16546 118832 16574
rect 121472 16546 122328 16574
rect 118804 480 118832 16546
rect 120632 14476 120684 14482
rect 120632 14418 120684 14424
rect 119896 6180 119948 6186
rect 119896 6122 119948 6128
rect 119908 480 119936 6122
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 14418
rect 122300 480 122328 16546
rect 123024 13116 123076 13122
rect 123024 13058 123076 13064
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 13058
rect 124680 3732 124732 3738
rect 124680 3674 124732 3680
rect 124692 480 124720 3674
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 156606
rect 133708 154465 133736 157383
rect 134628 156262 134656 158199
rect 135916 157010 135944 158471
rect 136086 157448 136142 157457
rect 136086 157383 136142 157392
rect 135904 157004 135956 157010
rect 135904 156946 135956 156952
rect 134616 156256 134668 156262
rect 134616 156198 134668 156204
rect 133694 154456 133750 154465
rect 133694 154391 133750 154400
rect 136100 154329 136128 157383
rect 137020 156942 137048 158471
rect 137008 156936 137060 156942
rect 137008 156878 137060 156884
rect 138400 156874 138428 158471
rect 138388 156868 138440 156874
rect 138388 156810 138440 156816
rect 139320 155961 139348 158607
rect 139674 158536 139730 158545
rect 139674 158471 139730 158480
rect 139688 156806 139716 158471
rect 141514 158264 141570 158273
rect 141514 158199 141570 158208
rect 141790 158264 141846 158273
rect 141790 158199 141846 158208
rect 146022 158264 146078 158273
rect 146022 158199 146078 158208
rect 146390 158264 146446 158273
rect 146390 158199 146446 158208
rect 150990 158264 151046 158273
rect 150990 158199 151046 158208
rect 140686 157992 140742 158001
rect 140686 157927 140742 157936
rect 139676 156800 139728 156806
rect 139676 156742 139728 156748
rect 139306 155952 139362 155961
rect 139306 155887 139362 155896
rect 140700 155582 140728 157927
rect 140688 155576 140740 155582
rect 140688 155518 140740 155524
rect 141528 154358 141556 158199
rect 141804 155786 141832 158199
rect 143078 157992 143134 158001
rect 143078 157927 143134 157936
rect 144550 157992 144606 158001
rect 144550 157927 144606 157936
rect 141792 155780 141844 155786
rect 141792 155722 141844 155728
rect 143092 155650 143120 157927
rect 143998 157448 144054 157457
rect 143998 157383 144054 157392
rect 143080 155644 143132 155650
rect 143080 155586 143132 155592
rect 144012 154834 144040 157383
rect 144564 155825 144592 157927
rect 145286 157720 145342 157729
rect 145286 157655 145342 157664
rect 144550 155816 144606 155825
rect 144550 155751 144606 155760
rect 145300 155446 145328 157655
rect 145288 155440 145340 155446
rect 145288 155382 145340 155388
rect 144000 154828 144052 154834
rect 144000 154770 144052 154776
rect 141516 154352 141568 154358
rect 136086 154320 136142 154329
rect 141516 154294 141568 154300
rect 136086 154255 136142 154264
rect 146036 154018 146064 158199
rect 146404 155378 146432 158199
rect 148690 158128 148746 158137
rect 148690 158063 148746 158072
rect 148414 157720 148470 157729
rect 148414 157655 148470 157664
rect 146392 155372 146444 155378
rect 146392 155314 146444 155320
rect 148428 155310 148456 157655
rect 148704 156126 148732 158063
rect 148782 157720 148838 157729
rect 148782 157655 148838 157664
rect 148692 156120 148744 156126
rect 148692 156062 148744 156068
rect 148796 155514 148824 157655
rect 149886 157448 149942 157457
rect 149886 157383 149942 157392
rect 148784 155508 148836 155514
rect 148784 155450 148836 155456
rect 148416 155304 148468 155310
rect 148416 155246 148468 155252
rect 149900 154290 149928 157383
rect 151004 155242 151032 158199
rect 159652 157962 159680 158607
rect 184018 158400 184074 158409
rect 184018 158335 184074 158344
rect 185950 158400 186006 158409
rect 185950 158335 186006 158344
rect 159640 157956 159692 157962
rect 159640 157898 159692 157904
rect 155774 157584 155830 157593
rect 155774 157519 155830 157528
rect 151358 157448 151414 157457
rect 151358 157383 151414 157392
rect 152646 157448 152702 157457
rect 152646 157383 152702 157392
rect 153842 157448 153898 157457
rect 153842 157383 153898 157392
rect 154486 157448 154542 157457
rect 154486 157383 154542 157392
rect 150992 155236 151044 155242
rect 150992 155178 151044 155184
rect 149888 154284 149940 154290
rect 149888 154226 149940 154232
rect 151372 154154 151400 157383
rect 151818 156632 151874 156641
rect 151818 156567 151874 156576
rect 151360 154148 151412 154154
rect 151360 154090 151412 154096
rect 146024 154012 146076 154018
rect 146024 153954 146076 153960
rect 129738 153776 129794 153785
rect 129738 153711 129794 153720
rect 128360 146940 128412 146946
rect 128360 146882 128412 146888
rect 126980 138712 127032 138718
rect 126980 138654 127032 138660
rect 126992 480 127020 138654
rect 127072 115252 127124 115258
rect 127072 115194 127124 115200
rect 127084 16574 127112 115194
rect 128372 16574 128400 146882
rect 129752 16574 129780 153711
rect 146300 151088 146352 151094
rect 146300 151030 146352 151036
rect 135260 148368 135312 148374
rect 135260 148310 135312 148316
rect 132500 142860 132552 142866
rect 132500 142802 132552 142808
rect 131120 127628 131172 127634
rect 131120 127570 131172 127576
rect 131132 16574 131160 127570
rect 132512 16574 132540 142802
rect 133880 122120 133932 122126
rect 133880 122062 133932 122068
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 122062
rect 135272 3806 135300 148310
rect 143540 144220 143592 144226
rect 143540 144162 143592 144168
rect 139400 141500 139452 141506
rect 139400 141442 139452 141448
rect 138020 126268 138072 126274
rect 138020 126210 138072 126216
rect 136640 120760 136692 120766
rect 136640 120702 136692 120708
rect 135352 101448 135404 101454
rect 135352 101390 135404 101396
rect 135260 3800 135312 3806
rect 135260 3742 135312 3748
rect 135364 3482 135392 101390
rect 136652 16574 136680 120702
rect 138032 16574 138060 126210
rect 139412 16574 139440 141442
rect 140780 119400 140832 119406
rect 140780 119342 140832 119348
rect 140792 16574 140820 119342
rect 142160 54528 142212 54534
rect 142160 54470 142212 54476
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 3800 136508 3806
rect 136456 3742 136508 3748
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3742
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 54470
rect 143552 480 143580 144162
rect 143632 116612 143684 116618
rect 143632 116554 143684 116560
rect 143644 16574 143672 116554
rect 144920 98660 144972 98666
rect 144920 98602 144972 98608
rect 144932 16574 144960 98602
rect 146312 16574 146340 151030
rect 150440 140140 150492 140146
rect 150440 140082 150492 140088
rect 147680 134564 147732 134570
rect 147680 134506 147732 134512
rect 147692 16574 147720 134506
rect 149060 129056 149112 129062
rect 149060 128998 149112 129004
rect 149072 16574 149100 128998
rect 150452 16574 150480 140082
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 9674 151860 156567
rect 152660 154426 152688 157383
rect 153856 154494 153884 157383
rect 153844 154488 153896 154494
rect 153844 154430 153896 154436
rect 152648 154420 152700 154426
rect 152648 154362 152700 154368
rect 154500 153610 154528 157383
rect 155788 154970 155816 157519
rect 157062 157448 157118 157457
rect 157062 157383 157118 157392
rect 155776 154964 155828 154970
rect 155776 154906 155828 154912
rect 157076 154086 157104 157383
rect 178038 156768 178094 156777
rect 178038 156703 178094 156712
rect 160098 155272 160154 155281
rect 160098 155207 160154 155216
rect 157064 154080 157116 154086
rect 157064 154022 157116 154028
rect 154488 153604 154540 153610
rect 154488 153546 154540 153552
rect 157340 149728 157392 149734
rect 157340 149670 157392 149676
rect 153200 145580 153252 145586
rect 153200 145522 153252 145528
rect 151912 117972 151964 117978
rect 151912 117914 151964 117920
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 117914
rect 153212 16574 153240 145522
rect 154580 144288 154632 144294
rect 154580 144230 154632 144236
rect 154592 16574 154620 144230
rect 155960 97300 156012 97306
rect 155960 97242 156012 97248
rect 155972 16574 156000 97242
rect 157352 16574 157380 149670
rect 158720 123480 158772 123486
rect 158720 123422 158772 123428
rect 158732 16574 158760 123422
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11830 160140 155207
rect 164240 153876 164292 153882
rect 164240 153818 164292 153824
rect 161480 137352 161532 137358
rect 161480 137294 161532 137300
rect 160192 17332 160244 17338
rect 160192 17274 160244 17280
rect 160100 11824 160152 11830
rect 160100 11766 160152 11772
rect 160204 6914 160232 17274
rect 161492 16574 161520 137294
rect 162860 113824 162912 113830
rect 162860 113766 162912 113772
rect 162872 16574 162900 113766
rect 164252 16574 164280 153818
rect 168380 152516 168432 152522
rect 168380 152458 168432 152464
rect 165620 135992 165672 135998
rect 165620 135934 165672 135940
rect 165632 16574 165660 135934
rect 167000 112464 167052 112470
rect 167000 112406 167052 112412
rect 167012 16574 167040 112406
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11824 161348 11830
rect 161296 11766 161348 11772
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11766
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 480 168420 152458
rect 175280 151156 175332 151162
rect 175280 151098 175332 151104
rect 168472 134632 168524 134638
rect 168472 134574 168524 134580
rect 168484 16574 168512 134574
rect 172520 133204 172572 133210
rect 172520 133146 172572 133152
rect 169760 124908 169812 124914
rect 169760 124850 169812 124856
rect 169772 16574 169800 124850
rect 172532 16574 172560 133146
rect 173900 111104 173952 111110
rect 173900 111046 173952 111052
rect 168484 16546 169616 16574
rect 169772 16546 170352 16574
rect 172532 16546 172744 16574
rect 169588 480 169616 16546
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171968 3800 172020 3806
rect 171968 3742 172020 3748
rect 171980 480 172008 3742
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 111046
rect 175292 16574 175320 151098
rect 176660 147008 176712 147014
rect 176660 146950 176712 146956
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 480 176700 146950
rect 178052 16574 178080 156703
rect 184032 156602 184060 158335
rect 184020 156596 184072 156602
rect 184020 156538 184072 156544
rect 185964 156534 185992 158335
rect 188724 157894 188752 158607
rect 191470 158264 191526 158273
rect 191470 158199 191526 158208
rect 195886 158264 195942 158273
rect 195886 158199 195942 158208
rect 188712 157888 188764 157894
rect 188712 157830 188764 157836
rect 185952 156528 186004 156534
rect 185952 156470 186004 156476
rect 191484 156466 191512 158199
rect 191472 156460 191524 156466
rect 191472 156402 191524 156408
rect 182178 155408 182234 155417
rect 182178 155343 182234 155352
rect 179420 131844 179472 131850
rect 179420 131786 179472 131792
rect 179432 16574 179460 131786
rect 180800 109744 180852 109750
rect 180800 109686 180852 109692
rect 180812 16574 180840 109686
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177856 15904 177908 15910
rect 177856 15846 177908 15852
rect 177868 480 177896 15846
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 155343
rect 195900 153950 195928 158199
rect 198462 157448 198518 157457
rect 198462 157383 198518 157392
rect 195888 153944 195940 153950
rect 195888 153886 195940 153892
rect 198476 153814 198504 157383
rect 198464 153808 198516 153814
rect 198464 153750 198516 153756
rect 193220 152584 193272 152590
rect 193220 152526 193272 152532
rect 184940 149796 184992 149802
rect 184940 149738 184992 149744
rect 183560 142928 183612 142934
rect 183560 142870 183612 142876
rect 183572 16574 183600 142870
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11830 184980 149738
rect 189080 148436 189132 148442
rect 189080 148378 189132 148384
rect 186320 130484 186372 130490
rect 186320 130426 186372 130432
rect 185032 108316 185084 108322
rect 185032 108258 185084 108264
rect 184940 11824 184992 11830
rect 184940 11766 184992 11772
rect 185044 6914 185072 108258
rect 186332 16574 186360 130426
rect 187700 105596 187752 105602
rect 187700 105538 187752 105544
rect 187712 16574 187740 105538
rect 189092 16574 189120 148378
rect 191840 133272 191892 133278
rect 191840 133214 191892 133220
rect 190460 129124 190512 129130
rect 190460 129066 190512 129072
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11766
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 129066
rect 191852 16574 191880 133214
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 152526
rect 195980 145648 196032 145654
rect 195980 145590 196032 145596
rect 193312 141568 193364 141574
rect 193312 141510 193364 141516
rect 193324 16574 193352 141510
rect 194600 53100 194652 53106
rect 194600 53042 194652 53048
rect 194612 16574 194640 53042
rect 195992 16574 196020 145590
rect 197360 140208 197412 140214
rect 197360 140150 197412 140156
rect 197372 16574 197400 140150
rect 198740 106956 198792 106962
rect 198740 106898 198792 106904
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 106898
rect 200132 16574 200160 159287
rect 206006 158672 206062 158681
rect 206006 158607 206062 158616
rect 206020 157826 206048 158607
rect 206008 157820 206060 157826
rect 206008 157762 206060 157768
rect 201038 157584 201094 157593
rect 201038 157519 201094 157528
rect 203430 157584 203486 157593
rect 203430 157519 203486 157528
rect 201052 155174 201080 157519
rect 201040 155168 201092 155174
rect 201040 155110 201092 155116
rect 203444 155106 203472 157519
rect 207018 156904 207074 156913
rect 207018 156839 207074 156848
rect 203432 155100 203484 155106
rect 203432 155042 203484 155048
rect 202880 153740 202932 153746
rect 202880 153682 202932 153688
rect 201500 138780 201552 138786
rect 201500 138722 201552 138728
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 138722
rect 201592 18624 201644 18630
rect 201592 18566 201644 18572
rect 201604 16574 201632 18566
rect 202892 16574 202920 153682
rect 204260 127696 204312 127702
rect 204260 127638 204312 127644
rect 204272 16574 204300 127638
rect 205640 104168 205692 104174
rect 205640 104110 205692 104116
rect 205652 16574 205680 104110
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 156839
rect 209780 151224 209832 151230
rect 209780 151166 209832 151172
rect 208400 126336 208452 126342
rect 208400 126278 208452 126284
rect 208412 16574 208440 126278
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 9674 209820 151166
rect 213920 149864 213972 149870
rect 213920 149806 213972 149812
rect 211160 137420 211212 137426
rect 211160 137362 211212 137368
rect 209872 19984 209924 19990
rect 209872 19926 209924 19932
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 19926
rect 211172 16574 211200 137362
rect 212540 21412 212592 21418
rect 212540 21354 212592 21360
rect 212552 16574 212580 21354
rect 213932 16574 213960 149806
rect 215300 148504 215352 148510
rect 215300 148446 215352 148452
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 148446
rect 219440 145716 219492 145722
rect 219440 145658 219492 145664
rect 218060 144356 218112 144362
rect 218060 144298 218112 144304
rect 216680 131912 216732 131918
rect 216680 131854 216732 131860
rect 216692 16574 216720 131854
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 144298
rect 218152 124976 218204 124982
rect 218152 124918 218204 124924
rect 218164 16574 218192 124918
rect 219452 16574 219480 145658
rect 220832 16574 220860 159326
rect 224958 155544 225014 155553
rect 224958 155479 225014 155488
rect 222200 136060 222252 136066
rect 222200 136002 222252 136008
rect 222212 16574 222240 136002
rect 223580 102876 223632 102882
rect 223580 102818 223632 102824
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 102818
rect 224972 16574 225000 155479
rect 229100 155032 229152 155038
rect 229100 154974 229152 154980
rect 227720 152652 227772 152658
rect 227720 152594 227772 152600
rect 226340 123548 226392 123554
rect 226340 123490 226392 123496
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 480 226380 123490
rect 227732 16574 227760 152594
rect 229112 16574 229140 154974
rect 231860 153672 231912 153678
rect 231860 153614 231912 153620
rect 230480 130552 230532 130558
rect 230480 130494 230532 130500
rect 230492 16574 230520 130494
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227536 4888 227588 4894
rect 227536 4830 227588 4836
rect 227548 480 227576 4830
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 153614
rect 233240 152720 233292 152726
rect 233240 152662 233292 152668
rect 233252 16574 233280 152662
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11830 234660 159394
rect 236000 142996 236052 143002
rect 236000 142938 236052 142944
rect 234712 100020 234764 100026
rect 234712 99962 234764 99968
rect 234620 11824 234672 11830
rect 234620 11766 234672 11772
rect 234724 6914 234752 99962
rect 236012 16574 236040 142938
rect 237760 32434 237788 306138
rect 237748 32428 237800 32434
rect 237748 32370 237800 32376
rect 236012 16546 236592 16574
rect 235816 11824 235868 11830
rect 235816 11766 235868 11772
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11766
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 238036 3738 238064 307022
rect 238128 159118 238156 307142
rect 238220 159225 238248 308343
rect 238312 306134 238340 310420
rect 238404 310406 238602 310434
rect 238404 306202 238432 310406
rect 238772 306542 238800 310420
rect 238970 310406 239076 310434
rect 238760 306536 238812 306542
rect 238760 306478 238812 306484
rect 239048 306354 239076 310406
rect 239128 306536 239180 306542
rect 239128 306478 239180 306484
rect 238956 306326 239076 306354
rect 238852 306264 238904 306270
rect 238852 306206 238904 306212
rect 238392 306196 238444 306202
rect 238392 306138 238444 306144
rect 238760 306196 238812 306202
rect 238760 306138 238812 306144
rect 238300 306128 238352 306134
rect 238300 306070 238352 306076
rect 238772 298790 238800 306138
rect 238864 300218 238892 306206
rect 238852 300212 238904 300218
rect 238852 300154 238904 300160
rect 238760 298784 238812 298790
rect 238760 298726 238812 298732
rect 238956 272542 238984 306326
rect 239036 306264 239088 306270
rect 239036 306206 239088 306212
rect 239048 293282 239076 306206
rect 239140 301578 239168 306478
rect 239128 301572 239180 301578
rect 239128 301514 239180 301520
rect 239036 293276 239088 293282
rect 239036 293218 239088 293224
rect 238944 272536 238996 272542
rect 238944 272478 238996 272484
rect 238300 267164 238352 267170
rect 238300 267106 238352 267112
rect 238206 159216 238262 159225
rect 238206 159151 238262 159160
rect 238116 159112 238168 159118
rect 238116 159054 238168 159060
rect 238312 158137 238340 267106
rect 238392 263084 238444 263090
rect 238392 263026 238444 263032
rect 238298 158128 238354 158137
rect 238298 158063 238354 158072
rect 238404 157826 238432 263026
rect 238484 250776 238536 250782
rect 238484 250718 238536 250724
rect 238496 157894 238524 250718
rect 238576 167680 238628 167686
rect 238576 167622 238628 167628
rect 238588 159730 238616 167622
rect 238576 159724 238628 159730
rect 238576 159666 238628 159672
rect 238484 157888 238536 157894
rect 238484 157830 238536 157836
rect 238392 157820 238444 157826
rect 238392 157762 238444 157768
rect 239232 89010 239260 310420
rect 239416 306474 239444 310420
rect 239404 306468 239456 306474
rect 239404 306410 239456 306416
rect 239600 306354 239628 310420
rect 239324 306326 239628 306354
rect 239692 310406 239890 310434
rect 239324 271182 239352 306326
rect 239692 306270 239720 310406
rect 239772 307828 239824 307834
rect 239772 307770 239824 307776
rect 239680 306264 239732 306270
rect 239680 306206 239732 306212
rect 239784 302234 239812 307770
rect 240060 306202 240088 310420
rect 240244 310406 240350 310434
rect 240048 306196 240100 306202
rect 240048 306138 240100 306144
rect 239416 302206 239812 302234
rect 239312 271176 239364 271182
rect 239312 271118 239364 271124
rect 239220 89004 239272 89010
rect 239220 88946 239272 88952
rect 239416 10334 239444 302206
rect 240244 269822 240272 310406
rect 240520 306354 240548 310420
rect 240704 307154 240732 310420
rect 240796 310406 240994 310434
rect 240692 307148 240744 307154
rect 240692 307090 240744 307096
rect 240796 306354 240824 310406
rect 240876 307896 240928 307902
rect 240876 307838 240928 307844
rect 240336 306326 240548 306354
rect 240704 306326 240824 306354
rect 240336 289202 240364 306326
rect 240416 306264 240468 306270
rect 240416 306206 240468 306212
rect 240428 297430 240456 306206
rect 240416 297424 240468 297430
rect 240416 297366 240468 297372
rect 240704 296714 240732 306326
rect 240888 302234 240916 307838
rect 241164 307834 241192 310420
rect 241152 307828 241204 307834
rect 241152 307770 241204 307776
rect 241348 306270 241376 310420
rect 241336 306264 241388 306270
rect 241336 306206 241388 306212
rect 240520 296686 240732 296714
rect 240796 302206 240916 302234
rect 240324 289196 240376 289202
rect 240324 289138 240376 289144
rect 240232 269816 240284 269822
rect 240232 269758 240284 269764
rect 240520 268394 240548 296686
rect 240508 268388 240560 268394
rect 240508 268330 240560 268336
rect 240796 159050 240824 302206
rect 241624 265674 241652 310420
rect 241808 307222 241836 310420
rect 241796 307216 241848 307222
rect 241796 307158 241848 307164
rect 241796 306400 241848 306406
rect 241992 306377 242020 310420
rect 242084 310406 242282 310434
rect 241796 306342 241848 306348
rect 241978 306368 242034 306377
rect 241704 306332 241756 306338
rect 241704 306274 241756 306280
rect 241716 283694 241744 306274
rect 241808 294710 241836 306342
rect 241978 306303 242034 306312
rect 241978 306096 242034 306105
rect 241978 306031 242034 306040
rect 241888 300484 241940 300490
rect 241888 300426 241940 300432
rect 241796 294704 241848 294710
rect 241796 294646 241848 294652
rect 241704 283688 241756 283694
rect 241704 283630 241756 283636
rect 241612 265668 241664 265674
rect 241612 265610 241664 265616
rect 241900 264246 241928 300426
rect 241992 296002 242020 306031
rect 242084 300490 242112 310406
rect 242256 308848 242308 308854
rect 242256 308790 242308 308796
rect 242164 307828 242216 307834
rect 242164 307770 242216 307776
rect 242072 300484 242124 300490
rect 242072 300426 242124 300432
rect 241980 295996 242032 296002
rect 241980 295938 242032 295944
rect 241888 264240 241940 264246
rect 241888 264182 241940 264188
rect 240784 159044 240836 159050
rect 240784 158986 240836 158992
rect 239404 10328 239456 10334
rect 239404 10270 239456 10276
rect 241704 9036 241756 9042
rect 241704 8978 241756 8984
rect 238116 6248 238168 6254
rect 238116 6190 238168 6196
rect 238024 3732 238076 3738
rect 238024 3674 238076 3680
rect 238128 480 238156 6190
rect 240508 4956 240560 4962
rect 240508 4898 240560 4904
rect 239312 3868 239364 3874
rect 239312 3810 239364 3816
rect 239324 480 239352 3810
rect 240520 480 240548 4898
rect 241716 480 241744 8978
rect 242176 7614 242204 307770
rect 242268 152522 242296 308790
rect 242452 306338 242480 310420
rect 242544 310406 242742 310434
rect 242544 306406 242572 310406
rect 242912 307834 242940 310420
rect 242900 307828 242952 307834
rect 242900 307770 242952 307776
rect 243096 306490 243124 310420
rect 243004 306462 243124 306490
rect 243188 310406 243386 310434
rect 242532 306400 242584 306406
rect 242532 306342 242584 306348
rect 242440 306332 242492 306338
rect 242440 306274 242492 306280
rect 243004 305658 243032 306462
rect 243188 306354 243216 310406
rect 243556 306354 243584 310420
rect 243740 308786 243768 310420
rect 243728 308780 243780 308786
rect 243728 308722 243780 308728
rect 243728 308644 243780 308650
rect 243728 308586 243780 308592
rect 243636 308100 243688 308106
rect 243636 308042 243688 308048
rect 243096 306326 243216 306354
rect 243280 306326 243584 306354
rect 242992 305652 243044 305658
rect 242992 305594 243044 305600
rect 243096 291922 243124 306326
rect 243176 306264 243228 306270
rect 243176 306206 243228 306212
rect 243084 291916 243136 291922
rect 243084 291858 243136 291864
rect 243188 261594 243216 306206
rect 243280 262954 243308 306326
rect 243648 305130 243676 308042
rect 243556 305102 243676 305130
rect 243268 262948 243320 262954
rect 243268 262890 243320 262896
rect 243176 261588 243228 261594
rect 243176 261530 243228 261536
rect 242256 152516 242308 152522
rect 242256 152458 242308 152464
rect 243556 8974 243584 305102
rect 243740 302234 243768 308586
rect 244016 305726 244044 310420
rect 244200 306270 244228 310420
rect 244188 306264 244240 306270
rect 244188 306206 244240 306212
rect 244004 305720 244056 305726
rect 244004 305662 244056 305668
rect 244384 304366 244412 310420
rect 244476 310406 244674 310434
rect 244372 304360 244424 304366
rect 244372 304302 244424 304308
rect 243648 302206 243768 302234
rect 243648 140078 243676 302206
rect 243636 140072 243688 140078
rect 243636 140014 243688 140020
rect 243544 8968 243596 8974
rect 243544 8910 243596 8916
rect 242164 7608 242216 7614
rect 242164 7550 242216 7556
rect 244096 3936 244148 3942
rect 244096 3878 244148 3884
rect 242900 3732 242952 3738
rect 242900 3674 242952 3680
rect 242912 480 242940 3674
rect 244108 480 244136 3878
rect 244476 3466 244504 310406
rect 244844 306354 244872 310420
rect 244568 306326 244872 306354
rect 244568 4826 244596 306326
rect 244740 306264 244792 306270
rect 244740 306206 244792 306212
rect 244648 10328 244700 10334
rect 244648 10270 244700 10276
rect 244556 4820 244608 4826
rect 244556 4762 244608 4768
rect 244660 3482 244688 10270
rect 244752 3602 244780 306206
rect 245120 303074 245148 310420
rect 245108 303068 245160 303074
rect 245108 303010 245160 303016
rect 245304 292574 245332 310420
rect 245488 306270 245516 310420
rect 245660 306536 245712 306542
rect 245660 306478 245712 306484
rect 245476 306264 245528 306270
rect 245476 306206 245528 306212
rect 245672 304434 245700 306478
rect 245660 304428 245712 304434
rect 245660 304370 245712 304376
rect 244844 292546 245332 292574
rect 244844 3602 244872 292546
rect 245764 280906 245792 310420
rect 245948 306542 245976 310420
rect 245936 306536 245988 306542
rect 245936 306478 245988 306484
rect 245844 306468 245896 306474
rect 245844 306410 245896 306416
rect 245856 286414 245884 306410
rect 246132 306354 246160 310420
rect 246408 308514 246436 310420
rect 246396 308508 246448 308514
rect 246396 308450 246448 308456
rect 246396 308032 246448 308038
rect 246396 307974 246448 307980
rect 246304 307896 246356 307902
rect 246304 307838 246356 307844
rect 245948 306326 246160 306354
rect 245948 297498 245976 306326
rect 246028 306264 246080 306270
rect 246028 306206 246080 306212
rect 245936 297492 245988 297498
rect 245936 297434 245988 297440
rect 245844 286408 245896 286414
rect 245844 286350 245896 286356
rect 245752 280900 245804 280906
rect 245752 280842 245804 280848
rect 246040 258806 246068 306206
rect 246028 258800 246080 258806
rect 246028 258742 246080 258748
rect 246316 22778 246344 307838
rect 246408 24138 246436 307974
rect 246592 306474 246620 310420
rect 246580 306468 246632 306474
rect 246580 306410 246632 306416
rect 246776 306270 246804 310420
rect 246856 307964 246908 307970
rect 246856 307906 246908 307912
rect 246764 306264 246816 306270
rect 246764 306206 246816 306212
rect 246868 292574 246896 307906
rect 247052 302234 247080 310420
rect 247236 303006 247264 310420
rect 247408 306400 247460 306406
rect 247408 306342 247460 306348
rect 247512 306354 247540 310420
rect 247696 308990 247724 310420
rect 247684 308984 247736 308990
rect 247684 308926 247736 308932
rect 247684 308508 247736 308514
rect 247684 308450 247736 308456
rect 247592 308168 247644 308174
rect 247592 308110 247644 308116
rect 247604 306490 247632 308110
rect 247696 307834 247724 308450
rect 247684 307828 247736 307834
rect 247684 307770 247736 307776
rect 247776 307828 247828 307834
rect 247776 307770 247828 307776
rect 247604 306462 247724 306490
rect 247316 306332 247368 306338
rect 247316 306274 247368 306280
rect 247224 303000 247276 303006
rect 247224 302942 247276 302948
rect 247052 302206 247264 302234
rect 246500 292546 246896 292574
rect 246500 137290 246528 292546
rect 247236 279546 247264 302206
rect 247328 285054 247356 306274
rect 247316 285048 247368 285054
rect 247316 284990 247368 284996
rect 247224 279540 247276 279546
rect 247224 279482 247276 279488
rect 246488 137284 246540 137290
rect 246488 137226 246540 137232
rect 247420 90370 247448 306342
rect 247512 306326 247632 306354
rect 247500 306264 247552 306270
rect 247500 306206 247552 306212
rect 247512 253298 247540 306206
rect 247604 296070 247632 306326
rect 247592 296064 247644 296070
rect 247592 296006 247644 296012
rect 247500 253292 247552 253298
rect 247500 253234 247552 253240
rect 247408 90364 247460 90370
rect 247408 90306 247460 90312
rect 246396 24132 246448 24138
rect 246396 24074 246448 24080
rect 246304 22772 246356 22778
rect 246304 22714 246356 22720
rect 247696 14482 247724 306462
rect 247788 130422 247816 307770
rect 247880 306338 247908 310420
rect 247972 310406 248170 310434
rect 247868 306332 247920 306338
rect 247868 306274 247920 306280
rect 247972 306270 248000 310406
rect 248340 306406 248368 310420
rect 248524 307834 248552 310420
rect 248512 307828 248564 307834
rect 248512 307770 248564 307776
rect 248328 306400 248380 306406
rect 248328 306342 248380 306348
rect 248512 306400 248564 306406
rect 248512 306342 248564 306348
rect 247960 306264 248012 306270
rect 247960 306206 248012 306212
rect 247776 130416 247828 130422
rect 247776 130358 247828 130364
rect 247684 14476 247736 14482
rect 247684 14418 247736 14424
rect 248524 11762 248552 306342
rect 248696 306332 248748 306338
rect 248696 306274 248748 306280
rect 248604 304156 248656 304162
rect 248604 304098 248656 304104
rect 248616 91798 248644 304098
rect 248708 135930 248736 306274
rect 248696 135924 248748 135930
rect 248696 135866 248748 135872
rect 248604 91792 248656 91798
rect 248604 91734 248656 91740
rect 248800 16574 248828 310420
rect 248984 307902 249012 310420
rect 249064 308576 249116 308582
rect 249064 308518 249116 308524
rect 248972 307896 249024 307902
rect 248972 307838 249024 307844
rect 249076 158982 249104 308518
rect 249168 306338 249196 310420
rect 249260 310406 249458 310434
rect 249260 306406 249288 310406
rect 249248 306400 249300 306406
rect 249248 306342 249300 306348
rect 249156 306332 249208 306338
rect 249156 306274 249208 306280
rect 249628 304162 249656 310420
rect 249904 307970 249932 310420
rect 250088 308106 250116 310420
rect 250076 308100 250128 308106
rect 250076 308042 250128 308048
rect 250272 308038 250300 310420
rect 250364 310406 250562 310434
rect 250260 308032 250312 308038
rect 250260 307974 250312 307980
rect 249892 307964 249944 307970
rect 249892 307906 249944 307912
rect 250364 306354 250392 310406
rect 250444 308236 250496 308242
rect 250444 308178 250496 308184
rect 249892 306332 249944 306338
rect 249892 306274 249944 306280
rect 249996 306326 250392 306354
rect 249616 304156 249668 304162
rect 249616 304098 249668 304104
rect 249064 158976 249116 158982
rect 249064 158918 249116 158924
rect 249904 94518 249932 306274
rect 249996 131782 250024 306326
rect 250076 306264 250128 306270
rect 250076 306206 250128 306212
rect 249984 131776 250036 131782
rect 249984 131718 250036 131724
rect 249892 94512 249944 94518
rect 249892 94454 249944 94460
rect 250088 86290 250116 306206
rect 250076 86284 250128 86290
rect 250076 86226 250128 86232
rect 248708 16546 248828 16574
rect 248512 11756 248564 11762
rect 248512 11698 248564 11704
rect 247592 7608 247644 7614
rect 247592 7550 247644 7556
rect 246396 4004 246448 4010
rect 246396 3946 246448 3952
rect 244740 3596 244792 3602
rect 244740 3538 244792 3544
rect 244832 3596 244884 3602
rect 244832 3538 244884 3544
rect 244464 3460 244516 3466
rect 244660 3454 245240 3482
rect 244464 3402 244516 3408
rect 245212 480 245240 3454
rect 246408 480 246436 3946
rect 247604 480 247632 7550
rect 248708 3670 248736 16546
rect 250456 13122 250484 308178
rect 250732 306338 250760 310420
rect 250720 306332 250772 306338
rect 250720 306274 250772 306280
rect 250916 306270 250944 310420
rect 250994 308680 251050 308689
rect 251192 308650 251220 310420
rect 250994 308615 251050 308624
rect 251180 308644 251232 308650
rect 250904 306264 250956 306270
rect 250904 306206 250956 306212
rect 251008 292574 251036 308615
rect 251180 308586 251232 308592
rect 251376 306762 251404 310420
rect 251192 306734 251404 306762
rect 251192 298654 251220 306734
rect 251560 306490 251588 310420
rect 251284 306462 251588 306490
rect 251652 310406 251850 310434
rect 251180 298648 251232 298654
rect 251180 298590 251232 298596
rect 250548 292546 251036 292574
rect 250548 158914 250576 292546
rect 250536 158908 250588 158914
rect 250536 158850 250588 158856
rect 251284 87650 251312 306462
rect 251652 306354 251680 310406
rect 251468 306326 251680 306354
rect 251364 298648 251416 298654
rect 251364 298590 251416 298596
rect 251376 93158 251404 298590
rect 251468 102814 251496 306326
rect 251548 304020 251600 304026
rect 251548 303962 251600 303968
rect 251560 141438 251588 303962
rect 252020 292574 252048 310420
rect 252296 308174 252324 310420
rect 252284 308168 252336 308174
rect 252284 308110 252336 308116
rect 252480 304026 252508 310420
rect 252664 308242 252692 310420
rect 252652 308236 252704 308242
rect 252652 308178 252704 308184
rect 252652 308100 252704 308106
rect 252652 308042 252704 308048
rect 252468 304020 252520 304026
rect 252468 303962 252520 303968
rect 251652 292546 252048 292574
rect 251548 141432 251600 141438
rect 251548 141374 251600 141380
rect 251456 102808 251508 102814
rect 251456 102750 251508 102756
rect 251364 93152 251416 93158
rect 251364 93094 251416 93100
rect 251272 87644 251324 87650
rect 251272 87586 251324 87592
rect 250444 13116 250496 13122
rect 250444 13058 250496 13064
rect 248788 7676 248840 7682
rect 248788 7618 248840 7624
rect 248696 3664 248748 3670
rect 248696 3606 248748 3612
rect 248800 480 248828 7618
rect 251652 6186 251680 292546
rect 252664 138718 252692 308042
rect 252940 307086 252968 310420
rect 252928 307080 252980 307086
rect 252928 307022 252980 307028
rect 253124 306354 253152 310420
rect 253308 308106 253336 310420
rect 253400 310406 253598 310434
rect 253296 308100 253348 308106
rect 253296 308042 253348 308048
rect 253400 307986 253428 310406
rect 253572 308644 253624 308650
rect 253572 308586 253624 308592
rect 252744 306332 252796 306338
rect 252744 306274 252796 306280
rect 252848 306326 253152 306354
rect 253216 307958 253428 307986
rect 252756 146946 252784 306274
rect 252848 156670 252876 306326
rect 253216 306218 253244 307958
rect 253388 307896 253440 307902
rect 253388 307838 253440 307844
rect 253296 307828 253348 307834
rect 253296 307770 253348 307776
rect 253124 306190 253244 306218
rect 253124 292574 253152 306190
rect 253308 292574 253336 307770
rect 252940 292546 253152 292574
rect 253216 292546 253336 292574
rect 252836 156664 252888 156670
rect 252836 156606 252888 156612
rect 252744 146940 252796 146946
rect 252744 146882 252796 146888
rect 252652 138712 252704 138718
rect 252652 138654 252704 138660
rect 252940 115258 252968 292546
rect 253216 142866 253244 292546
rect 253296 156664 253348 156670
rect 253296 156606 253348 156612
rect 253204 142860 253256 142866
rect 253204 142802 253256 142808
rect 252928 115252 252980 115258
rect 252928 115194 252980 115200
rect 251640 6180 251692 6186
rect 251640 6122 251692 6128
rect 253308 4010 253336 156606
rect 253400 155281 253428 307838
rect 253584 307834 253612 308586
rect 253572 307828 253624 307834
rect 253572 307770 253624 307776
rect 253768 306338 253796 310420
rect 253966 310406 254072 310434
rect 253756 306332 253808 306338
rect 253756 306274 253808 306280
rect 254044 304842 254072 310406
rect 254136 310406 254242 310434
rect 254032 304836 254084 304842
rect 254032 304778 254084 304784
rect 254032 304700 254084 304706
rect 254032 304642 254084 304648
rect 253386 155272 253442 155281
rect 253386 155207 253442 155216
rect 253388 146940 253440 146946
rect 253388 146882 253440 146888
rect 253296 4004 253348 4010
rect 253296 3946 253348 3952
rect 253400 3874 253428 146882
rect 254044 122126 254072 304642
rect 254136 127634 254164 310406
rect 254412 308650 254440 310420
rect 254504 310406 254702 310434
rect 254400 308644 254452 308650
rect 254400 308586 254452 308592
rect 254216 306332 254268 306338
rect 254216 306274 254268 306280
rect 254228 148374 254256 306274
rect 254308 304836 254360 304842
rect 254308 304778 254360 304784
rect 254320 153785 254348 304778
rect 254504 304706 254532 310406
rect 254492 304700 254544 304706
rect 254492 304642 254544 304648
rect 254872 302234 254900 310420
rect 254952 307828 255004 307834
rect 254952 307770 255004 307776
rect 254412 302206 254900 302234
rect 254306 153776 254362 153785
rect 254306 153711 254362 153720
rect 254216 148368 254268 148374
rect 254216 148310 254268 148316
rect 254124 127628 254176 127634
rect 254124 127570 254176 127576
rect 254032 122120 254084 122126
rect 254032 122062 254084 122068
rect 254412 101454 254440 302206
rect 254964 296714 254992 307770
rect 255056 306338 255084 310420
rect 255044 306332 255096 306338
rect 255044 306274 255096 306280
rect 255332 306218 255360 310420
rect 255516 306320 255544 310420
rect 255700 307834 255728 310420
rect 255688 307828 255740 307834
rect 255688 307770 255740 307776
rect 255780 306332 255832 306338
rect 255516 306292 255728 306320
rect 255332 306190 255636 306218
rect 255504 306128 255556 306134
rect 255504 306070 255556 306076
rect 255412 306060 255464 306066
rect 255412 306002 255464 306008
rect 254596 296686 254992 296714
rect 254596 141506 254624 296686
rect 254584 141500 254636 141506
rect 254584 141442 254636 141448
rect 254584 122120 254636 122126
rect 254584 122062 254636 122068
rect 254400 101448 254452 101454
rect 254400 101390 254452 101396
rect 254596 3942 254624 122062
rect 255424 116618 255452 306002
rect 255516 119406 255544 306070
rect 255608 120766 255636 306190
rect 255700 126274 255728 306292
rect 255780 306274 255832 306280
rect 255792 144226 255820 306274
rect 255976 306134 256004 310420
rect 255964 306128 256016 306134
rect 255964 306070 256016 306076
rect 256160 305980 256188 310420
rect 256240 307828 256292 307834
rect 256240 307770 256292 307776
rect 255884 305952 256188 305980
rect 255780 144220 255832 144226
rect 255780 144162 255832 144168
rect 255688 126268 255740 126274
rect 255688 126210 255740 126216
rect 255596 120760 255648 120766
rect 255596 120702 255648 120708
rect 255504 119400 255556 119406
rect 255504 119342 255556 119348
rect 255412 116612 255464 116618
rect 255412 116554 255464 116560
rect 255884 54534 255912 305952
rect 256252 302234 256280 307770
rect 256344 306338 256372 310420
rect 256436 310406 256634 310434
rect 256332 306332 256384 306338
rect 256332 306274 256384 306280
rect 256436 306066 256464 310406
rect 256804 306320 256832 310420
rect 257080 307018 257108 310420
rect 257068 307012 257120 307018
rect 257068 306954 257120 306960
rect 257160 306808 257212 306814
rect 257160 306750 257212 306756
rect 256712 306292 256832 306320
rect 256884 306332 256936 306338
rect 256424 306060 256476 306066
rect 256424 306002 256476 306008
rect 255976 302206 256280 302234
rect 255976 145586 256004 302206
rect 255964 145580 256016 145586
rect 255964 145522 256016 145528
rect 256712 98666 256740 306292
rect 256884 306274 256936 306280
rect 256792 306128 256844 306134
rect 256792 306070 256844 306076
rect 256804 117978 256832 306070
rect 256896 129062 256924 306274
rect 257068 306196 257120 306202
rect 257068 306138 257120 306144
rect 256976 304292 257028 304298
rect 256976 304234 257028 304240
rect 256988 134570 257016 304234
rect 257080 140146 257108 306138
rect 257172 151094 257200 306750
rect 257264 304298 257292 310420
rect 257344 308712 257396 308718
rect 257344 308654 257396 308660
rect 257252 304292 257304 304298
rect 257252 304234 257304 304240
rect 257160 151088 257212 151094
rect 257160 151030 257212 151036
rect 257068 140140 257120 140146
rect 257068 140082 257120 140088
rect 256976 134564 257028 134570
rect 256976 134506 257028 134512
rect 256884 129056 256936 129062
rect 256884 128998 256936 129004
rect 256792 117972 256844 117978
rect 256792 117914 256844 117920
rect 256700 98660 256752 98666
rect 256700 98602 256752 98608
rect 255872 54528 255924 54534
rect 255872 54470 255924 54476
rect 257356 12510 257384 308654
rect 257448 306338 257476 310420
rect 257540 310406 257738 310434
rect 257436 306332 257488 306338
rect 257436 306274 257488 306280
rect 257540 306202 257568 310406
rect 257528 306196 257580 306202
rect 257528 306138 257580 306144
rect 257908 306134 257936 310420
rect 258106 310406 258304 310434
rect 258276 306490 258304 310406
rect 258368 307834 258396 310420
rect 258356 307828 258408 307834
rect 258356 307770 258408 307776
rect 258276 306462 258488 306490
rect 258172 306332 258224 306338
rect 258172 306274 258224 306280
rect 257896 306128 257948 306134
rect 257896 306070 257948 306076
rect 258184 123486 258212 306274
rect 258356 306196 258408 306202
rect 258356 306138 258408 306144
rect 258264 302660 258316 302666
rect 258264 302602 258316 302608
rect 258276 144294 258304 302602
rect 258368 149734 258396 306138
rect 258460 156641 258488 306462
rect 258552 302666 258580 310420
rect 258540 302660 258592 302666
rect 258540 302602 258592 302608
rect 258736 296714 258764 310420
rect 258828 310406 259026 310434
rect 258828 306202 258856 310406
rect 259196 306338 259224 310420
rect 259184 306332 259236 306338
rect 259184 306274 259236 306280
rect 259472 306202 259500 310420
rect 259656 307902 259684 310420
rect 259644 307896 259696 307902
rect 259644 307838 259696 307844
rect 259840 306746 259868 310420
rect 259932 310406 260130 310434
rect 259828 306740 259880 306746
rect 259828 306682 259880 306688
rect 259932 306626 259960 310406
rect 260300 307986 260328 310420
rect 259656 306598 259960 306626
rect 260024 307958 260328 307986
rect 259552 306400 259604 306406
rect 259552 306342 259604 306348
rect 258816 306196 258868 306202
rect 258816 306138 258868 306144
rect 259460 306196 259512 306202
rect 259460 306138 259512 306144
rect 258552 296686 258764 296714
rect 258446 156632 258502 156641
rect 258446 156567 258502 156576
rect 258356 149728 258408 149734
rect 258356 149670 258408 149676
rect 258264 144288 258316 144294
rect 258264 144230 258316 144236
rect 258172 123480 258224 123486
rect 258172 123422 258224 123428
rect 258552 97306 258580 296686
rect 259564 112470 259592 306342
rect 259656 113830 259684 306598
rect 259828 306468 259880 306474
rect 259828 306410 259880 306416
rect 259736 306332 259788 306338
rect 259736 306274 259788 306280
rect 259748 135998 259776 306274
rect 259840 137358 259868 306410
rect 260024 306320 260052 307958
rect 260104 307896 260156 307902
rect 260104 307838 260156 307844
rect 259932 306292 260052 306320
rect 259932 153882 259960 306292
rect 260012 306196 260064 306202
rect 260012 306138 260064 306144
rect 259920 153876 259972 153882
rect 259920 153818 259972 153824
rect 259828 137352 259880 137358
rect 259828 137294 259880 137300
rect 259736 135992 259788 135998
rect 259736 135934 259788 135940
rect 259644 113824 259696 113830
rect 259644 113766 259696 113772
rect 259552 112464 259604 112470
rect 259552 112406 259604 112412
rect 258540 97300 258592 97306
rect 258540 97242 258592 97248
rect 260024 17338 260052 306138
rect 260116 156777 260144 307838
rect 260484 306338 260512 310420
rect 260576 310406 260774 310434
rect 260576 306406 260604 310406
rect 260944 308854 260972 310420
rect 260932 308848 260984 308854
rect 260932 308790 260984 308796
rect 260564 306400 260616 306406
rect 260564 306342 260616 306348
rect 260472 306332 260524 306338
rect 260472 306274 260524 306280
rect 260932 305244 260984 305250
rect 260932 305186 260984 305192
rect 260102 156768 260158 156777
rect 260102 156703 260158 156712
rect 260102 141400 260158 141409
rect 260102 141335 260158 141344
rect 260012 17332 260064 17338
rect 260012 17274 260064 17280
rect 259552 17264 259604 17270
rect 259552 17206 259604 17212
rect 259564 16574 259592 17206
rect 259564 16546 260052 16574
rect 255872 12504 255924 12510
rect 255872 12446 255924 12452
rect 257344 12504 257396 12510
rect 257344 12446 257396 12452
rect 254676 6180 254728 6186
rect 254676 6122 254728 6128
rect 254584 3936 254636 3942
rect 254584 3878 254636 3884
rect 253388 3868 253440 3874
rect 253388 3810 253440 3816
rect 251180 3664 251232 3670
rect 251180 3606 251232 3612
rect 249984 3596 250036 3602
rect 249984 3538 250036 3544
rect 249996 480 250024 3538
rect 251192 480 251220 3606
rect 253480 3528 253532 3534
rect 253480 3470 253532 3476
rect 252376 3460 252428 3466
rect 252376 3402 252428 3408
rect 252388 480 252416 3402
rect 253492 480 253520 3470
rect 254688 480 254716 6122
rect 255884 480 255912 12446
rect 257068 4140 257120 4146
rect 257068 4082 257120 4088
rect 257080 480 257108 4082
rect 258172 3868 258224 3874
rect 258172 3810 258224 3816
rect 258184 3602 258212 3810
rect 258172 3596 258224 3602
rect 258172 3538 258224 3544
rect 258264 3596 258316 3602
rect 258264 3538 258316 3544
rect 258276 480 258304 3538
rect 260024 3482 260052 16546
rect 260116 3602 260144 141335
rect 260944 111110 260972 305186
rect 261036 124914 261064 310490
rect 261142 310406 261340 310434
rect 261208 307964 261260 307970
rect 261208 307906 261260 307912
rect 261116 177336 261168 177342
rect 261116 177278 261168 177284
rect 261024 124908 261076 124914
rect 261024 124850 261076 124856
rect 260932 111104 260984 111110
rect 260932 111046 260984 111052
rect 261128 16574 261156 177278
rect 261220 133210 261248 307906
rect 261312 134638 261340 310406
rect 261588 306320 261616 310420
rect 261680 310406 261878 310434
rect 261680 307970 261708 310406
rect 261668 307964 261720 307970
rect 261668 307906 261720 307912
rect 261668 307828 261720 307834
rect 261668 307770 261720 307776
rect 261404 306292 261616 306320
rect 261300 134632 261352 134638
rect 261300 134574 261352 134580
rect 261208 133204 261260 133210
rect 261208 133146 261260 133152
rect 261128 16546 261340 16574
rect 260196 13184 260248 13190
rect 260196 13126 260248 13132
rect 260208 4146 260236 13126
rect 260196 4140 260248 4146
rect 260196 4082 260248 4088
rect 260104 3596 260156 3602
rect 260104 3538 260156 3544
rect 261312 3482 261340 16546
rect 261404 3806 261432 306292
rect 261680 302234 261708 307770
rect 262048 305250 262076 310420
rect 262232 307834 262260 310420
rect 262220 307828 262272 307834
rect 262220 307770 262272 307776
rect 262404 306400 262456 306406
rect 262404 306342 262456 306348
rect 262312 306264 262364 306270
rect 262312 306206 262364 306212
rect 262036 305244 262088 305250
rect 262036 305186 262088 305192
rect 261496 302206 261708 302234
rect 261496 151162 261524 302206
rect 261484 151156 261536 151162
rect 261484 151098 261536 151104
rect 261484 133204 261536 133210
rect 261484 133146 261536 133152
rect 261392 3800 261444 3806
rect 261392 3742 261444 3748
rect 261496 3670 261524 133146
rect 262324 109750 262352 306206
rect 262416 131850 262444 306342
rect 262508 147014 262536 310420
rect 262588 306332 262640 306338
rect 262588 306274 262640 306280
rect 262600 155417 262628 306274
rect 262586 155408 262642 155417
rect 262586 155343 262642 155352
rect 262496 147008 262548 147014
rect 262496 146950 262548 146956
rect 262404 131844 262456 131850
rect 262404 131786 262456 131792
rect 262312 109744 262364 109750
rect 262312 109686 262364 109692
rect 262692 15910 262720 310420
rect 262876 307902 262904 310420
rect 262968 310406 263166 310434
rect 262864 307896 262916 307902
rect 262864 307838 262916 307844
rect 262968 306406 262996 310406
rect 262956 306400 263008 306406
rect 262956 306342 263008 306348
rect 263336 306270 263364 310420
rect 263520 306338 263548 310420
rect 263508 306332 263560 306338
rect 263508 306274 263560 306280
rect 263692 306332 263744 306338
rect 263692 306274 263744 306280
rect 263324 306264 263376 306270
rect 263324 306206 263376 306212
rect 263600 302796 263652 302802
rect 263600 302738 263652 302744
rect 263612 105602 263640 302738
rect 263704 108322 263732 306274
rect 263796 306082 263824 310420
rect 263980 306338 264008 310420
rect 264072 310406 264270 310434
rect 263968 306332 264020 306338
rect 263968 306274 264020 306280
rect 263968 306128 264020 306134
rect 263796 306054 263916 306082
rect 263968 306070 264020 306076
rect 263784 305992 263836 305998
rect 263784 305934 263836 305940
rect 263796 130490 263824 305934
rect 263888 142934 263916 306054
rect 263980 148442 264008 306070
rect 264072 149802 264100 310406
rect 264244 307080 264296 307086
rect 264244 307022 264296 307028
rect 264060 149796 264112 149802
rect 264060 149738 264112 149744
rect 263968 148436 264020 148442
rect 263968 148378 264020 148384
rect 263876 142928 263928 142934
rect 263876 142870 263928 142876
rect 263784 130484 263836 130490
rect 263784 130426 263836 130432
rect 263692 108316 263744 108322
rect 263692 108258 263744 108264
rect 263600 105596 263652 105602
rect 263600 105538 263652 105544
rect 262680 15904 262732 15910
rect 262680 15846 262732 15852
rect 264152 14476 264204 14482
rect 264152 14418 264204 14424
rect 261484 3664 261536 3670
rect 261484 3606 261536 3612
rect 260024 3454 260696 3482
rect 261312 3454 261800 3482
rect 259460 3324 259512 3330
rect 259460 3266 259512 3272
rect 259472 480 259500 3266
rect 260668 480 260696 3454
rect 261772 480 261800 3454
rect 262956 3392 263008 3398
rect 262956 3334 263008 3340
rect 262968 480 262996 3334
rect 264164 480 264192 14418
rect 264256 3738 264284 307022
rect 264440 305998 264468 310420
rect 264428 305992 264480 305998
rect 264428 305934 264480 305940
rect 264624 302802 264652 310420
rect 264716 310406 264914 310434
rect 264716 306134 264744 310406
rect 264704 306128 264756 306134
rect 264704 306070 264756 306076
rect 264980 303476 265032 303482
rect 264980 303418 265032 303424
rect 264612 302796 264664 302802
rect 264612 302738 264664 302744
rect 264334 148336 264390 148345
rect 264334 148271 264390 148280
rect 264244 3732 264296 3738
rect 264244 3674 264296 3680
rect 264348 3330 264376 148271
rect 264992 53106 265020 303418
rect 265084 129130 265112 310420
rect 265268 306354 265296 310420
rect 265176 306326 265296 306354
rect 265452 310406 265558 310434
rect 265348 306332 265400 306338
rect 265176 133278 265204 306326
rect 265348 306274 265400 306280
rect 265256 306264 265308 306270
rect 265256 306206 265308 306212
rect 265268 141574 265296 306206
rect 265360 145654 265388 306274
rect 265452 152590 265480 310406
rect 265624 307828 265676 307834
rect 265624 307770 265676 307776
rect 265636 159361 265664 307770
rect 265728 306270 265756 310420
rect 265716 306264 265768 306270
rect 265716 306206 265768 306212
rect 265912 303482 265940 310420
rect 266004 310406 266202 310434
rect 266464 310406 266662 310434
rect 266004 306338 266032 310406
rect 265992 306332 266044 306338
rect 265992 306274 266044 306280
rect 265900 303476 265952 303482
rect 265900 303418 265952 303424
rect 265622 159352 265678 159361
rect 265622 159287 265678 159296
rect 265440 152584 265492 152590
rect 265440 152526 265492 152532
rect 265348 145648 265400 145654
rect 265348 145590 265400 145596
rect 265624 145580 265676 145586
rect 265624 145522 265676 145528
rect 265256 141568 265308 141574
rect 265256 141510 265308 141516
rect 265164 133272 265216 133278
rect 265164 133214 265216 133220
rect 265072 129124 265124 129130
rect 265072 129066 265124 129072
rect 265162 129024 265218 129033
rect 265162 128959 265218 128968
rect 264980 53100 265032 53106
rect 264980 53042 265032 53048
rect 264336 3324 264388 3330
rect 264336 3266 264388 3272
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265176 354 265204 128959
rect 265636 3874 265664 145522
rect 266464 106962 266492 310406
rect 266636 306332 266688 306338
rect 266636 306274 266688 306280
rect 266544 306264 266596 306270
rect 266544 306206 266596 306212
rect 266556 127702 266584 306206
rect 266648 138786 266676 306274
rect 266740 140214 266768 310490
rect 266832 307834 266860 310420
rect 266820 307828 266872 307834
rect 266820 307770 266872 307776
rect 266820 306400 266872 306406
rect 266820 306342 266872 306348
rect 266832 153746 266860 306342
rect 267016 306338 267044 310420
rect 267108 310406 267306 310434
rect 267004 306332 267056 306338
rect 267004 306274 267056 306280
rect 267108 292574 267136 310406
rect 267476 306406 267504 310420
rect 267464 306400 267516 306406
rect 267464 306342 267516 306348
rect 267660 306270 267688 310420
rect 267844 310406 267950 310434
rect 267740 306400 267792 306406
rect 267740 306342 267792 306348
rect 267648 306264 267700 306270
rect 267648 306206 267700 306212
rect 266924 292546 267136 292574
rect 266820 153740 266872 153746
rect 266820 153682 266872 153688
rect 266728 140208 266780 140214
rect 266728 140150 266780 140156
rect 266636 138780 266688 138786
rect 266636 138722 266688 138728
rect 266544 127696 266596 127702
rect 266544 127638 266596 127644
rect 266452 106956 266504 106962
rect 266452 106898 266504 106904
rect 266924 18630 266952 292546
rect 267752 19990 267780 306342
rect 267844 104174 267872 310406
rect 268120 307018 268148 310420
rect 268108 307012 268160 307018
rect 268108 306954 268160 306960
rect 268200 306808 268252 306814
rect 268200 306750 268252 306756
rect 268016 306332 268068 306338
rect 268016 306274 268068 306280
rect 267924 300552 267976 300558
rect 267924 300494 267976 300500
rect 267936 126342 267964 300494
rect 268028 137426 268056 306274
rect 268108 306264 268160 306270
rect 268108 306206 268160 306212
rect 268120 151230 268148 306206
rect 268212 156913 268240 306750
rect 268304 300558 268332 310420
rect 268396 310406 268594 310434
rect 268396 306406 268424 310406
rect 268476 307896 268528 307902
rect 268476 307838 268528 307844
rect 268384 306400 268436 306406
rect 268384 306342 268436 306348
rect 268292 300552 268344 300558
rect 268292 300494 268344 300500
rect 268488 292574 268516 307838
rect 268764 306270 268792 310420
rect 268856 310406 269054 310434
rect 268856 306338 268884 310406
rect 269224 306354 269252 310420
rect 269422 310406 269620 310434
rect 268844 306332 268896 306338
rect 268844 306274 268896 306280
rect 269132 306326 269252 306354
rect 269396 306400 269448 306406
rect 269396 306342 269448 306348
rect 269304 306332 269356 306338
rect 268752 306264 268804 306270
rect 268752 306206 268804 306212
rect 268396 292546 268516 292574
rect 268198 156904 268254 156913
rect 268198 156839 268254 156848
rect 268108 151224 268160 151230
rect 268108 151166 268160 151172
rect 268200 150476 268252 150482
rect 268200 150418 268252 150424
rect 268016 137420 268068 137426
rect 268016 137362 268068 137368
rect 267924 126336 267976 126342
rect 267924 126278 267976 126284
rect 267832 104168 267884 104174
rect 267832 104110 267884 104116
rect 267740 19984 267792 19990
rect 267740 19926 267792 19932
rect 266912 18624 266964 18630
rect 266912 18566 266964 18572
rect 266544 11756 266596 11762
rect 266544 11698 266596 11704
rect 265624 3868 265676 3874
rect 265624 3810 265676 3816
rect 266556 480 266584 11698
rect 268212 6914 268240 150418
rect 268396 7682 268424 292546
rect 269132 21418 269160 306326
rect 269304 306274 269356 306280
rect 269212 306264 269264 306270
rect 269212 306206 269264 306212
rect 269224 124982 269252 306206
rect 269316 131918 269344 306274
rect 269408 144362 269436 306342
rect 269592 297498 269620 310406
rect 269580 297492 269632 297498
rect 269580 297434 269632 297440
rect 269580 297288 269632 297294
rect 269580 297230 269632 297236
rect 269488 291168 269540 291174
rect 269488 291110 269540 291116
rect 269500 148510 269528 291110
rect 269592 149870 269620 297230
rect 269684 291174 269712 310420
rect 269764 307828 269816 307834
rect 269764 307770 269816 307776
rect 269672 291168 269724 291174
rect 269672 291110 269724 291116
rect 269776 152658 269804 307770
rect 269868 306338 269896 310420
rect 270052 306406 270080 310420
rect 270144 310406 270342 310434
rect 270040 306400 270092 306406
rect 270040 306342 270092 306348
rect 269856 306332 269908 306338
rect 269856 306274 269908 306280
rect 270144 306270 270172 310406
rect 270132 306264 270184 306270
rect 270132 306206 270184 306212
rect 270512 306105 270540 310420
rect 270696 306270 270724 310420
rect 270788 310406 270986 310434
rect 270684 306264 270736 306270
rect 270684 306206 270736 306212
rect 270498 306096 270554 306105
rect 270498 306031 270554 306040
rect 270592 305992 270644 305998
rect 270592 305934 270644 305940
rect 270500 305856 270552 305862
rect 270500 305798 270552 305804
rect 269856 303408 269908 303414
rect 269856 303350 269908 303356
rect 269868 154018 269896 303350
rect 269948 303272 270000 303278
rect 269948 303214 270000 303220
rect 269960 155310 269988 303214
rect 270040 303204 270092 303210
rect 270040 303146 270092 303152
rect 269948 155304 270000 155310
rect 269948 155246 270000 155252
rect 270052 155242 270080 303146
rect 270040 155236 270092 155242
rect 270040 155178 270092 155184
rect 269856 154012 269908 154018
rect 269856 153954 269908 153960
rect 269764 152652 269816 152658
rect 269764 152594 269816 152600
rect 269580 149864 269632 149870
rect 269580 149806 269632 149812
rect 269488 148504 269540 148510
rect 269488 148446 269540 148452
rect 269396 144356 269448 144362
rect 269396 144298 269448 144304
rect 269764 144084 269816 144090
rect 269764 144026 269816 144032
rect 269304 131912 269356 131918
rect 269304 131854 269356 131860
rect 269212 124976 269264 124982
rect 269212 124918 269264 124924
rect 269120 21412 269172 21418
rect 269120 21354 269172 21360
rect 268384 7676 268436 7682
rect 268384 7618 268436 7624
rect 268212 6886 268424 6914
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 267752 480 267780 3538
rect 265318 354 265430 480
rect 265176 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 6886
rect 269776 3534 269804 144026
rect 269856 124908 269908 124914
rect 269856 124850 269908 124856
rect 269764 3528 269816 3534
rect 269764 3470 269816 3476
rect 269868 3398 269896 124850
rect 270512 4894 270540 305798
rect 270604 102882 270632 305934
rect 270684 305924 270736 305930
rect 270684 305866 270736 305872
rect 270696 123554 270724 305866
rect 270788 136066 270816 310406
rect 271156 306490 271184 310420
rect 270880 306462 271184 306490
rect 271248 310406 271446 310434
rect 270880 306202 270908 306462
rect 271248 306354 271276 310406
rect 270972 306326 271276 306354
rect 270868 306196 270920 306202
rect 270868 306138 270920 306144
rect 270866 306096 270922 306105
rect 270866 306031 270922 306040
rect 270880 145722 270908 306031
rect 270972 155553 271000 306326
rect 271052 306264 271104 306270
rect 271052 306206 271104 306212
rect 271064 159390 271092 306206
rect 271616 305930 271644 310420
rect 271604 305924 271656 305930
rect 271604 305866 271656 305872
rect 271800 305862 271828 310420
rect 272076 307834 272104 310420
rect 272064 307828 272116 307834
rect 272064 307770 272116 307776
rect 272064 306468 272116 306474
rect 272064 306410 272116 306416
rect 271972 306332 272024 306338
rect 271972 306274 272024 306280
rect 271788 305856 271840 305862
rect 271788 305798 271840 305804
rect 271052 159384 271104 159390
rect 271052 159326 271104 159332
rect 271144 155916 271196 155922
rect 271144 155858 271196 155864
rect 270958 155544 271014 155553
rect 270958 155479 271014 155488
rect 270868 145716 270920 145722
rect 270868 145658 270920 145664
rect 270776 136060 270828 136066
rect 270776 136002 270828 136008
rect 270684 123548 270736 123554
rect 270684 123490 270736 123496
rect 270592 102876 270644 102882
rect 270592 102818 270644 102824
rect 270500 4888 270552 4894
rect 270500 4830 270552 4836
rect 271156 3466 271184 155858
rect 271984 130558 272012 306274
rect 272076 152726 272104 306410
rect 272156 306400 272208 306406
rect 272156 306342 272208 306348
rect 272168 153678 272196 306342
rect 272260 155038 272288 310420
rect 272444 306338 272472 310420
rect 272536 310406 272734 310434
rect 272536 306406 272564 310406
rect 272904 306474 272932 310420
rect 272892 306468 272944 306474
rect 272892 306410 272944 306416
rect 272524 306400 272576 306406
rect 273088 306354 273116 310420
rect 272524 306342 272576 306348
rect 272432 306332 272484 306338
rect 272432 306274 272484 306280
rect 272628 306326 273116 306354
rect 273260 306332 273312 306338
rect 272628 306218 272656 306326
rect 273260 306274 273312 306280
rect 272352 306190 272656 306218
rect 272248 155032 272300 155038
rect 272248 154974 272300 154980
rect 272156 153672 272208 153678
rect 272156 153614 272208 153620
rect 272064 152720 272116 152726
rect 272064 152662 272116 152668
rect 271972 130552 272024 130558
rect 271972 130494 272024 130500
rect 272352 100026 272380 306190
rect 272524 303544 272576 303550
rect 272524 303486 272576 303492
rect 272536 154358 272564 303486
rect 272800 303476 272852 303482
rect 272800 303418 272852 303424
rect 272614 303104 272670 303113
rect 272614 303039 272670 303048
rect 272628 155961 272656 303039
rect 272614 155952 272670 155961
rect 272614 155887 272670 155896
rect 272812 155825 272840 303418
rect 272798 155816 272854 155825
rect 272798 155751 272854 155760
rect 272524 154352 272576 154358
rect 272524 154294 272576 154300
rect 272524 151836 272576 151842
rect 272524 151778 272576 151784
rect 272340 100020 272392 100026
rect 272340 99962 272392 99968
rect 272432 10532 272484 10538
rect 272432 10474 272484 10480
rect 271236 8288 271288 8294
rect 271236 8230 271288 8236
rect 271144 3460 271196 3466
rect 271144 3402 271196 3408
rect 269856 3392 269908 3398
rect 269856 3334 269908 3340
rect 270040 3052 270092 3058
rect 270040 2994 270092 3000
rect 270052 480 270080 2994
rect 271248 480 271276 8230
rect 272444 480 272472 10474
rect 272536 3058 272564 151778
rect 273272 4962 273300 306274
rect 273364 306270 273392 310420
rect 273444 306468 273496 306474
rect 273444 306410 273496 306416
rect 273352 306264 273404 306270
rect 273352 306206 273404 306212
rect 273456 306082 273484 306410
rect 273364 306054 273484 306082
rect 273364 6254 273392 306054
rect 273444 304020 273496 304026
rect 273444 303962 273496 303968
rect 273456 9042 273484 303962
rect 273548 143002 273576 310420
rect 273640 310406 273838 310434
rect 273640 306474 273668 310406
rect 273628 306468 273680 306474
rect 273628 306410 273680 306416
rect 274008 306354 274036 310420
rect 274088 307964 274140 307970
rect 274088 307906 274140 307912
rect 273640 306326 274036 306354
rect 273640 146946 273668 306326
rect 273720 306264 273772 306270
rect 273720 306206 273772 306212
rect 273732 159458 273760 306206
rect 274100 302234 274128 307906
rect 274192 306338 274220 310420
rect 274284 310406 274482 310434
rect 274180 306332 274232 306338
rect 274180 306274 274232 306280
rect 274284 304026 274312 310406
rect 274652 307086 274680 310420
rect 274640 307080 274692 307086
rect 274640 307022 274692 307028
rect 274732 306332 274784 306338
rect 274732 306274 274784 306280
rect 274272 304020 274324 304026
rect 274272 303962 274324 303968
rect 273916 302206 274128 302234
rect 273720 159452 273772 159458
rect 273720 159394 273772 159400
rect 273916 150482 273944 302206
rect 273904 150476 273956 150482
rect 273904 150418 273956 150424
rect 273902 147656 273958 147665
rect 273902 147591 273958 147600
rect 273628 146940 273680 146946
rect 273628 146882 273680 146888
rect 273536 142996 273588 143002
rect 273536 142938 273588 142944
rect 273444 9036 273496 9042
rect 273444 8978 273496 8984
rect 273352 6248 273404 6254
rect 273352 6190 273404 6196
rect 273260 4956 273312 4962
rect 273260 4898 273312 4904
rect 273916 3602 273944 147591
rect 274744 10334 274772 306274
rect 274836 122126 274864 310420
rect 274928 310406 275126 310434
rect 274928 306338 274956 310406
rect 275296 306354 275324 310420
rect 274916 306332 274968 306338
rect 274916 306274 274968 306280
rect 275020 306326 275324 306354
rect 274916 306196 274968 306202
rect 274916 306138 274968 306144
rect 274928 145586 274956 306138
rect 275020 156670 275048 306326
rect 275480 305572 275508 310420
rect 275560 308780 275612 308786
rect 275560 308722 275612 308728
rect 275112 305544 275508 305572
rect 275008 156664 275060 156670
rect 275008 156606 275060 156612
rect 274916 145580 274968 145586
rect 274916 145522 274968 145528
rect 275008 145580 275060 145586
rect 275008 145522 275060 145528
rect 274824 122120 274876 122126
rect 274824 122062 274876 122068
rect 274732 10328 274784 10334
rect 274732 10270 274784 10276
rect 273904 3596 273956 3602
rect 273904 3538 273956 3544
rect 273628 3120 273680 3126
rect 273628 3062 273680 3068
rect 272524 3052 272576 3058
rect 272524 2994 272576 3000
rect 273640 480 273668 3062
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 354 274906 480
rect 275020 354 275048 145522
rect 275112 7614 275140 305544
rect 275572 305402 275600 308722
rect 275756 307902 275784 310420
rect 275744 307896 275796 307902
rect 275744 307838 275796 307844
rect 275940 306202 275968 310420
rect 276138 310406 276244 310434
rect 275928 306196 275980 306202
rect 275928 306138 275980 306144
rect 275296 305374 275600 305402
rect 275296 8294 275324 305374
rect 275928 303612 275980 303618
rect 275928 303554 275980 303560
rect 275376 303000 275428 303006
rect 275376 302942 275428 302948
rect 275388 155174 275416 302942
rect 275468 302932 275520 302938
rect 275468 302874 275520 302880
rect 275376 155168 275428 155174
rect 275376 155110 275428 155116
rect 275480 155106 275508 302874
rect 275836 297696 275888 297702
rect 275836 297638 275888 297644
rect 275848 158030 275876 297638
rect 275940 158166 275968 303554
rect 276112 303068 276164 303074
rect 276112 303010 276164 303016
rect 276020 158704 276072 158710
rect 276020 158646 276072 158652
rect 276032 158409 276060 158646
rect 276018 158400 276074 158409
rect 276018 158335 276074 158344
rect 275928 158160 275980 158166
rect 275928 158102 275980 158108
rect 275836 158024 275888 158030
rect 275836 157966 275888 157972
rect 276020 155848 276072 155854
rect 276020 155790 276072 155796
rect 276032 155378 276060 155790
rect 276020 155372 276072 155378
rect 276020 155314 276072 155320
rect 275468 155100 275520 155106
rect 275468 155042 275520 155048
rect 276020 154556 276072 154562
rect 276020 154498 276072 154504
rect 276032 154222 276060 154498
rect 276020 154216 276072 154222
rect 276020 154158 276072 154164
rect 276124 13190 276152 303010
rect 276216 133210 276244 310406
rect 276400 309134 276428 310420
rect 276400 309106 276520 309134
rect 276296 304292 276348 304298
rect 276296 304234 276348 304240
rect 276308 144090 276336 304234
rect 276492 299474 276520 309106
rect 276584 304298 276612 310420
rect 276676 310406 276874 310434
rect 276572 304292 276624 304298
rect 276572 304234 276624 304240
rect 276400 299446 276520 299474
rect 276400 155922 276428 299446
rect 276676 296714 276704 310406
rect 277044 308718 277072 310420
rect 277032 308712 277084 308718
rect 277032 308654 277084 308660
rect 276940 306196 276992 306202
rect 276940 306138 276992 306144
rect 276952 302234 276980 306138
rect 277032 306128 277084 306134
rect 277032 306070 277084 306076
rect 277044 302682 277072 306070
rect 277124 306060 277176 306066
rect 277124 306002 277176 306008
rect 277136 302870 277164 306002
rect 277228 303074 277256 310420
rect 277504 308009 277532 310420
rect 277490 308000 277546 308009
rect 277490 307935 277546 307944
rect 277688 307873 277716 310420
rect 277674 307864 277730 307873
rect 277674 307799 277730 307808
rect 277872 306354 277900 310420
rect 277400 306332 277452 306338
rect 277400 306274 277452 306280
rect 277504 306326 277900 306354
rect 277964 310406 278162 310434
rect 277308 305720 277360 305726
rect 277308 305662 277360 305668
rect 277216 303068 277268 303074
rect 277216 303010 277268 303016
rect 277320 302954 277348 305662
rect 277228 302926 277348 302954
rect 277124 302864 277176 302870
rect 277124 302806 277176 302812
rect 277044 302654 277164 302682
rect 276952 302206 277072 302234
rect 276492 296686 276704 296714
rect 276388 155916 276440 155922
rect 276388 155858 276440 155864
rect 276296 144084 276348 144090
rect 276296 144026 276348 144032
rect 276204 133204 276256 133210
rect 276204 133146 276256 133152
rect 276112 13184 276164 13190
rect 276112 13126 276164 13132
rect 276020 13116 276072 13122
rect 276020 13058 276072 13064
rect 275284 8288 275336 8294
rect 275284 8230 275336 8236
rect 275100 7608 275152 7614
rect 275100 7550 275152 7556
rect 276032 480 276060 13058
rect 276492 6186 276520 296686
rect 277044 161474 277072 302206
rect 276860 161446 277072 161474
rect 276860 158642 276888 161446
rect 276572 158636 276624 158642
rect 276572 158578 276624 158584
rect 276848 158636 276900 158642
rect 276848 158578 276900 158584
rect 276584 158137 276612 158578
rect 277136 158409 277164 302654
rect 277122 158400 277178 158409
rect 277122 158335 277178 158344
rect 276570 158128 276626 158137
rect 276570 158063 276626 158072
rect 277228 155854 277256 302926
rect 277308 302864 277360 302870
rect 277308 302806 277360 302812
rect 277216 155848 277268 155854
rect 277216 155790 277268 155796
rect 277320 154222 277348 302806
rect 277308 154216 277360 154222
rect 277308 154158 277360 154164
rect 277412 14482 277440 306274
rect 277504 17270 277532 306326
rect 277584 306264 277636 306270
rect 277584 306206 277636 306212
rect 277596 124914 277624 306206
rect 277964 296714 277992 310406
rect 278044 307828 278096 307834
rect 278044 307770 278096 307776
rect 277688 296686 277992 296714
rect 277688 177342 277716 296686
rect 277676 177336 277728 177342
rect 277676 177278 277728 177284
rect 277584 124908 277636 124914
rect 277584 124850 277636 124856
rect 277492 17264 277544 17270
rect 277492 17206 277544 17212
rect 277400 14476 277452 14482
rect 277400 14418 277452 14424
rect 278056 11762 278084 307770
rect 278332 306270 278360 310420
rect 278516 306338 278544 310420
rect 278792 307873 278820 310420
rect 278872 307896 278924 307902
rect 278778 307864 278834 307873
rect 278872 307838 278924 307844
rect 278778 307799 278834 307808
rect 278504 306332 278556 306338
rect 278504 306274 278556 306280
rect 278320 306264 278372 306270
rect 278320 306206 278372 306212
rect 278320 305652 278372 305658
rect 278320 305594 278372 305600
rect 278136 303136 278188 303142
rect 278136 303078 278188 303084
rect 278148 153950 278176 303078
rect 278228 303068 278280 303074
rect 278228 303010 278280 303016
rect 278136 153944 278188 153950
rect 278136 153886 278188 153892
rect 278240 153814 278268 303010
rect 278332 158273 278360 305594
rect 278884 302234 278912 307838
rect 278976 307834 279004 310420
rect 279252 307873 279280 310420
rect 279436 307970 279464 310420
rect 279424 307964 279476 307970
rect 279424 307906 279476 307912
rect 279238 307864 279294 307873
rect 278964 307828 279016 307834
rect 279238 307799 279294 307808
rect 278964 307770 279016 307776
rect 279620 306354 279648 310420
rect 279896 308786 279924 310420
rect 279884 308780 279936 308786
rect 279884 308722 279936 308728
rect 279884 308644 279936 308650
rect 279884 308586 279936 308592
rect 279792 307964 279844 307970
rect 279792 307906 279844 307912
rect 279700 307828 279752 307834
rect 279700 307770 279752 307776
rect 278792 302206 278912 302234
rect 278976 306326 279648 306354
rect 278686 300248 278742 300257
rect 278686 300183 278742 300192
rect 278596 297832 278648 297838
rect 278596 297774 278648 297780
rect 278318 158264 278374 158273
rect 278318 158199 278374 158208
rect 278608 157078 278636 297774
rect 278700 158545 278728 300183
rect 278686 158536 278742 158545
rect 278686 158471 278742 158480
rect 278596 157072 278648 157078
rect 278596 157014 278648 157020
rect 278228 153808 278280 153814
rect 278228 153750 278280 153756
rect 278136 124500 278188 124506
rect 278136 124442 278188 124448
rect 278044 11756 278096 11762
rect 278044 11698 278096 11704
rect 276480 6180 276532 6186
rect 276480 6122 276532 6128
rect 277124 4140 277176 4146
rect 277124 4082 277176 4088
rect 277136 480 277164 4082
rect 278148 3126 278176 124442
rect 278792 16574 278820 302206
rect 278976 151842 279004 306326
rect 279330 306232 279386 306241
rect 279330 306167 279386 306176
rect 278964 151836 279016 151842
rect 278964 151778 279016 151784
rect 278792 16546 279096 16574
rect 278320 4208 278372 4214
rect 278320 4150 278372 4156
rect 278136 3120 278188 3126
rect 278136 3062 278188 3068
rect 278332 480 278360 4150
rect 274794 326 275048 354
rect 274794 -960 274906 326
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 279344 10538 279372 306167
rect 279712 302234 279740 307770
rect 279804 305130 279832 307906
rect 279896 305402 279924 308586
rect 280080 306241 280108 310420
rect 280066 306232 280122 306241
rect 280066 306167 280122 306176
rect 279896 305374 280108 305402
rect 279804 305102 280016 305130
rect 279884 303340 279936 303346
rect 279884 303282 279936 303288
rect 279436 302206 279740 302234
rect 279332 10532 279384 10538
rect 279332 10474 279384 10480
rect 279436 4214 279464 302206
rect 279698 300656 279754 300665
rect 279698 300591 279754 300600
rect 279608 300212 279660 300218
rect 279608 300154 279660 300160
rect 279620 155582 279648 300154
rect 279608 155576 279660 155582
rect 279608 155518 279660 155524
rect 279712 155446 279740 300591
rect 279790 300384 279846 300393
rect 279790 300319 279846 300328
rect 279700 155440 279752 155446
rect 279700 155382 279752 155388
rect 279804 154562 279832 300319
rect 279792 154556 279844 154562
rect 279792 154498 279844 154504
rect 279896 154290 279924 303282
rect 279988 156874 280016 305102
rect 280080 157146 280108 305374
rect 280068 157140 280120 157146
rect 280068 157082 280120 157088
rect 279976 156868 280028 156874
rect 279976 156810 280028 156816
rect 279988 156398 280016 156810
rect 280080 156806 280108 157082
rect 280068 156800 280120 156806
rect 280068 156742 280120 156748
rect 279976 156392 280028 156398
rect 279976 156334 280028 156340
rect 280068 154556 280120 154562
rect 280068 154498 280120 154504
rect 279884 154284 279936 154290
rect 279884 154226 279936 154232
rect 280080 154154 280108 154498
rect 280068 154148 280120 154154
rect 280068 154090 280120 154096
rect 279516 146600 279568 146606
rect 279516 146542 279568 146548
rect 279424 4208 279476 4214
rect 279424 4150 279476 4156
rect 279528 4146 279556 146542
rect 280264 124506 280292 310420
rect 280356 310406 280554 310434
rect 280356 145586 280384 310406
rect 280436 306332 280488 306338
rect 280436 306274 280488 306280
rect 280448 146606 280476 306274
rect 280724 296714 280752 310420
rect 280908 306338 280936 310420
rect 281184 307834 281212 310420
rect 281368 307902 281396 310420
rect 281448 308236 281500 308242
rect 281448 308178 281500 308184
rect 281356 307896 281408 307902
rect 281356 307838 281408 307844
rect 281172 307828 281224 307834
rect 281172 307770 281224 307776
rect 280896 306332 280948 306338
rect 280896 306274 280948 306280
rect 280988 306332 281040 306338
rect 280988 306274 281040 306280
rect 281000 306134 281028 306274
rect 280988 306128 281040 306134
rect 280988 306070 281040 306076
rect 281080 305992 281132 305998
rect 281080 305934 281132 305940
rect 280988 305924 281040 305930
rect 280988 305866 281040 305872
rect 280896 305856 280948 305862
rect 280896 305798 280948 305804
rect 280804 305788 280856 305794
rect 280804 305730 280856 305736
rect 280540 296686 280752 296714
rect 280436 146600 280488 146606
rect 280436 146542 280488 146548
rect 280344 145580 280396 145586
rect 280344 145522 280396 145528
rect 280344 125588 280396 125594
rect 280344 125530 280396 125536
rect 280252 124500 280304 124506
rect 280252 124442 280304 124448
rect 280356 6914 280384 125530
rect 280540 13122 280568 296686
rect 280816 156466 280844 305730
rect 280908 156534 280936 305798
rect 281000 156602 281028 305866
rect 281092 157321 281120 305934
rect 281354 300520 281410 300529
rect 281354 300455 281410 300464
rect 281078 157312 281134 157321
rect 281078 157247 281134 157256
rect 280988 156596 281040 156602
rect 280988 156538 281040 156544
rect 280896 156528 280948 156534
rect 280896 156470 280948 156476
rect 280804 156460 280856 156466
rect 280804 156402 280856 156408
rect 281368 154358 281396 300455
rect 281356 154352 281408 154358
rect 281356 154294 281408 154300
rect 280528 13116 280580 13122
rect 280528 13058 280580 13064
rect 280356 6886 280752 6914
rect 279516 4140 279568 4146
rect 279516 4082 279568 4088
rect 280724 480 280752 6886
rect 281460 3602 281488 308178
rect 281644 306474 281672 310420
rect 281828 306626 281856 310420
rect 281736 306598 281856 306626
rect 281632 306468 281684 306474
rect 281632 306410 281684 306416
rect 281736 306354 281764 306598
rect 281552 306326 281764 306354
rect 281448 3596 281500 3602
rect 281448 3538 281500 3544
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 306326
rect 282012 306218 282040 310420
rect 281644 306190 282040 306218
rect 282104 310406 282302 310434
rect 281644 3534 281672 306190
rect 281724 306128 281776 306134
rect 282104 306082 282132 310406
rect 282184 306468 282236 306474
rect 282184 306410 282236 306416
rect 281724 306070 281776 306076
rect 281736 4214 281764 306070
rect 281828 306054 282132 306082
rect 281828 5574 281856 306054
rect 282196 305946 282224 306410
rect 282472 306134 282500 310420
rect 282656 308378 282684 310420
rect 282828 308916 282880 308922
rect 282828 308858 282880 308864
rect 282644 308372 282696 308378
rect 282644 308314 282696 308320
rect 282460 306128 282512 306134
rect 282460 306070 282512 306076
rect 282736 306128 282788 306134
rect 282736 306070 282788 306076
rect 282644 306060 282696 306066
rect 282644 306002 282696 306008
rect 281920 305918 282224 305946
rect 281920 125594 281948 305918
rect 282552 300416 282604 300422
rect 282552 300358 282604 300364
rect 282460 297764 282512 297770
rect 282460 297706 282512 297712
rect 282472 158438 282500 297706
rect 282460 158432 282512 158438
rect 282460 158374 282512 158380
rect 282564 157214 282592 300358
rect 282552 157208 282604 157214
rect 282552 157150 282604 157156
rect 282656 155718 282684 306002
rect 282368 155712 282420 155718
rect 282368 155654 282420 155660
rect 282644 155712 282696 155718
rect 282644 155654 282696 155660
rect 282380 155514 282408 155654
rect 282748 155650 282776 306070
rect 282840 157010 282868 308858
rect 282932 306218 282960 310420
rect 283116 306354 283144 310420
rect 283314 310406 283512 310434
rect 283116 306326 283328 306354
rect 282932 306190 283236 306218
rect 283012 305584 283064 305590
rect 283012 305526 283064 305532
rect 282828 157004 282880 157010
rect 282828 156946 282880 156952
rect 282920 156732 282972 156738
rect 282920 156674 282972 156680
rect 282932 156194 282960 156674
rect 282920 156188 282972 156194
rect 282920 156130 282972 156136
rect 282736 155644 282788 155650
rect 282736 155586 282788 155592
rect 282368 155508 282420 155514
rect 282368 155450 282420 155456
rect 282920 155508 282972 155514
rect 282920 155450 282972 155456
rect 282932 154834 282960 155450
rect 282920 154828 282972 154834
rect 282920 154770 282972 154776
rect 281908 125588 281960 125594
rect 281908 125530 281960 125536
rect 283024 6798 283052 305526
rect 283208 299474 283236 306190
rect 283116 299446 283236 299474
rect 283116 294794 283144 299446
rect 283116 294766 283236 294794
rect 283104 294636 283156 294642
rect 283104 294578 283156 294584
rect 283116 6934 283144 294578
rect 283208 145586 283236 294766
rect 283300 294642 283328 306326
rect 283288 294636 283340 294642
rect 283288 294578 283340 294584
rect 283196 145580 283248 145586
rect 283196 145522 283248 145528
rect 283104 6928 283156 6934
rect 283104 6870 283156 6876
rect 283012 6792 283064 6798
rect 283012 6734 283064 6740
rect 281816 5568 281868 5574
rect 281816 5510 281868 5516
rect 283484 4962 283512 310406
rect 283576 308038 283604 310420
rect 283656 308372 283708 308378
rect 283656 308314 283708 308320
rect 283564 308032 283616 308038
rect 283564 307974 283616 307980
rect 283668 292574 283696 308314
rect 283760 308242 283788 310420
rect 283932 308848 283984 308854
rect 283932 308790 283984 308796
rect 283748 308236 283800 308242
rect 283748 308178 283800 308184
rect 283748 308100 283800 308106
rect 283748 308042 283800 308048
rect 283760 303090 283788 308042
rect 283944 305454 283972 308790
rect 284036 307834 284064 310420
rect 284116 309120 284168 309126
rect 284116 309062 284168 309068
rect 284024 307828 284076 307834
rect 284024 307770 284076 307776
rect 283932 305448 283984 305454
rect 283932 305390 283984 305396
rect 284128 303634 284156 309062
rect 284220 305590 284248 310420
rect 284404 308106 284432 310420
rect 284392 308100 284444 308106
rect 284392 308042 284444 308048
rect 284680 307902 284708 310420
rect 284668 307896 284720 307902
rect 284668 307838 284720 307844
rect 284864 306354 284892 310420
rect 284944 307828 284996 307834
rect 284944 307770 284996 307776
rect 284312 306326 284892 306354
rect 284208 305584 284260 305590
rect 284208 305526 284260 305532
rect 284208 305448 284260 305454
rect 284208 305390 284260 305396
rect 284036 303606 284156 303634
rect 284036 303362 284064 303606
rect 284036 303334 284156 303362
rect 283760 303062 284064 303090
rect 283840 300484 283892 300490
rect 283840 300426 283892 300432
rect 283576 292546 283696 292574
rect 283576 155922 283604 292546
rect 283852 158273 283880 300426
rect 283932 297628 283984 297634
rect 283932 297570 283984 297576
rect 283838 158264 283894 158273
rect 283838 158199 283894 158208
rect 283852 158098 283880 158199
rect 283840 158092 283892 158098
rect 283840 158034 283892 158040
rect 283748 157344 283800 157350
rect 283748 157286 283800 157292
rect 283760 156874 283788 157286
rect 283748 156868 283800 156874
rect 283748 156810 283800 156816
rect 283564 155916 283616 155922
rect 283564 155858 283616 155864
rect 283944 154086 283972 297570
rect 284036 157350 284064 303062
rect 284024 157344 284076 157350
rect 284024 157286 284076 157292
rect 284128 156738 284156 303334
rect 284116 156732 284168 156738
rect 284116 156674 284168 156680
rect 284220 155514 284248 305390
rect 284208 155508 284260 155514
rect 284208 155450 284260 155456
rect 283932 154080 283984 154086
rect 283932 154022 283984 154028
rect 284208 5568 284260 5574
rect 284208 5510 284260 5516
rect 283472 4956 283524 4962
rect 283472 4898 283524 4904
rect 281724 4208 281776 4214
rect 281724 4150 281776 4156
rect 281632 3528 281684 3534
rect 281632 3470 281684 3476
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 284220 3482 284248 5510
rect 284312 4826 284340 306326
rect 284392 305584 284444 305590
rect 284392 305526 284444 305532
rect 284404 151230 284432 305526
rect 284484 305516 284536 305522
rect 284484 305458 284536 305464
rect 284496 159662 284524 305458
rect 284484 159656 284536 159662
rect 284484 159598 284536 159604
rect 284484 157344 284536 157350
rect 284484 157286 284536 157292
rect 284496 156126 284524 157286
rect 284484 156120 284536 156126
rect 284484 156062 284536 156068
rect 284392 151224 284444 151230
rect 284392 151166 284444 151172
rect 284956 11830 284984 307770
rect 285048 305522 285076 310420
rect 285140 310406 285338 310434
rect 285140 305590 285168 310406
rect 285220 308032 285272 308038
rect 285220 307974 285272 307980
rect 285128 305584 285180 305590
rect 285128 305526 285180 305532
rect 285036 305516 285088 305522
rect 285036 305458 285088 305464
rect 285232 302234 285260 307974
rect 285508 307873 285536 310420
rect 285706 310406 285904 310434
rect 285588 308780 285640 308786
rect 285588 308722 285640 308728
rect 285494 307864 285550 307873
rect 285494 307799 285550 307808
rect 285048 302206 285260 302234
rect 285048 140214 285076 302206
rect 285220 300824 285272 300830
rect 285220 300766 285272 300772
rect 285232 171086 285260 300766
rect 285404 300756 285456 300762
rect 285404 300698 285456 300704
rect 285312 300144 285364 300150
rect 285312 300086 285364 300092
rect 285220 171080 285272 171086
rect 285220 171022 285272 171028
rect 285232 170406 285260 171022
rect 285220 170400 285272 170406
rect 285220 170342 285272 170348
rect 285324 161474 285352 300086
rect 285140 161446 285352 161474
rect 285140 157962 285168 161446
rect 285128 157956 285180 157962
rect 285128 157898 285180 157904
rect 285140 157593 285168 157898
rect 285126 157584 285182 157593
rect 285126 157519 285182 157528
rect 285416 157282 285444 300698
rect 285496 300348 285548 300354
rect 285496 300290 285548 300296
rect 285404 157276 285456 157282
rect 285404 157218 285456 157224
rect 285508 155786 285536 300290
rect 285600 157350 285628 308722
rect 285876 306626 285904 310406
rect 285968 306762 285996 310420
rect 285968 306734 286088 306762
rect 285876 306598 285996 306626
rect 285680 306468 285732 306474
rect 285680 306410 285732 306416
rect 285588 157344 285640 157350
rect 285588 157286 285640 157292
rect 285496 155780 285548 155786
rect 285496 155722 285548 155728
rect 285036 140208 285088 140214
rect 285036 140150 285088 140156
rect 285692 13122 285720 306410
rect 285772 306400 285824 306406
rect 285772 306342 285824 306348
rect 285784 141506 285812 306342
rect 285968 302234 285996 306598
rect 285876 302206 285996 302234
rect 285876 297498 285904 302206
rect 285864 297492 285916 297498
rect 285864 297434 285916 297440
rect 286060 297378 286088 306734
rect 286152 306406 286180 310420
rect 286244 310406 286442 310434
rect 286140 306400 286192 306406
rect 286140 306342 286192 306348
rect 285876 297350 286088 297378
rect 285876 149870 285904 297350
rect 285956 297288 286008 297294
rect 285956 297230 286008 297236
rect 285968 156534 285996 297230
rect 286244 292574 286272 310406
rect 286416 308984 286468 308990
rect 286416 308926 286468 308932
rect 286324 307896 286376 307902
rect 286324 307838 286376 307844
rect 286060 292546 286272 292574
rect 285956 156528 286008 156534
rect 285956 156470 286008 156476
rect 285956 155916 286008 155922
rect 285956 155858 286008 155864
rect 285864 149864 285916 149870
rect 285864 149806 285916 149812
rect 285772 141500 285824 141506
rect 285772 141442 285824 141448
rect 285968 16574 285996 155858
rect 286060 155174 286088 292546
rect 286140 158092 286192 158098
rect 286140 158034 286192 158040
rect 286152 157758 286180 158034
rect 286140 157752 286192 157758
rect 286140 157694 286192 157700
rect 286140 156936 286192 156942
rect 286140 156878 286192 156884
rect 286152 156262 286180 156878
rect 286140 156256 286192 156262
rect 286140 156198 286192 156204
rect 286140 155916 286192 155922
rect 286140 155858 286192 155864
rect 286152 155446 286180 155858
rect 286140 155440 286192 155446
rect 286140 155382 286192 155388
rect 286048 155168 286100 155174
rect 286048 155110 286100 155116
rect 285968 16546 286272 16574
rect 285680 13116 285732 13122
rect 285680 13058 285732 13064
rect 284944 11824 284996 11830
rect 284944 11766 284996 11772
rect 284300 4820 284352 4826
rect 284300 4762 284352 4768
rect 285404 4208 285456 4214
rect 285404 4150 285456 4156
rect 283116 480 283144 3470
rect 284220 3454 284340 3482
rect 284312 480 284340 3454
rect 285416 480 285444 4150
rect 286244 3482 286272 16546
rect 286336 4894 286364 307838
rect 286428 158846 286456 308926
rect 286612 306474 286640 310420
rect 286796 307834 286824 310420
rect 286784 307828 286836 307834
rect 286784 307770 286836 307776
rect 287072 306474 287100 310420
rect 287256 307018 287284 310420
rect 287244 307012 287296 307018
rect 287244 306954 287296 306960
rect 287336 306808 287388 306814
rect 287336 306750 287388 306756
rect 287152 306536 287204 306542
rect 287152 306478 287204 306484
rect 286600 306468 286652 306474
rect 286600 306410 286652 306416
rect 287060 306468 287112 306474
rect 287060 306410 287112 306416
rect 287060 305516 287112 305522
rect 287060 305458 287112 305464
rect 286968 300620 287020 300626
rect 286968 300562 287020 300568
rect 286876 300076 286928 300082
rect 286876 300018 286928 300024
rect 286692 248192 286744 248198
rect 286692 248134 286744 248140
rect 286704 238754 286732 248134
rect 286784 247444 286836 247450
rect 286784 247386 286836 247392
rect 286796 247081 286824 247386
rect 286782 247072 286838 247081
rect 286782 247007 286838 247016
rect 286704 238726 286824 238754
rect 286796 159186 286824 238726
rect 286784 159180 286836 159186
rect 286784 159122 286836 159128
rect 286416 158840 286468 158846
rect 286416 158782 286468 158788
rect 286888 158098 286916 300018
rect 286876 158092 286928 158098
rect 286876 158034 286928 158040
rect 286980 156942 287008 300562
rect 286968 156936 287020 156942
rect 286968 156878 287020 156884
rect 287072 11762 287100 305458
rect 287164 14482 287192 306478
rect 287244 305584 287296 305590
rect 287244 305526 287296 305532
rect 287256 145722 287284 305526
rect 287348 147014 287376 306750
rect 287440 306542 287468 310420
rect 287532 310406 287730 310434
rect 287428 306536 287480 306542
rect 287428 306478 287480 306484
rect 287428 306400 287480 306406
rect 287428 306342 287480 306348
rect 287440 153882 287468 306342
rect 287532 156602 287560 310406
rect 287704 308712 287756 308718
rect 287704 308654 287756 308660
rect 287716 307970 287744 308654
rect 287704 307964 287756 307970
rect 287704 307906 287756 307912
rect 287612 306468 287664 306474
rect 287612 306410 287664 306416
rect 287624 159594 287652 306410
rect 287900 305590 287928 310420
rect 287888 305584 287940 305590
rect 287888 305526 287940 305532
rect 288084 305522 288112 310420
rect 288176 310406 288374 310434
rect 288558 310406 288664 310434
rect 288176 306406 288204 310406
rect 288532 306468 288584 306474
rect 288532 306410 288584 306416
rect 288164 306400 288216 306406
rect 288164 306342 288216 306348
rect 288440 306400 288492 306406
rect 288440 306342 288492 306348
rect 288072 305516 288124 305522
rect 288072 305458 288124 305464
rect 288256 300008 288308 300014
rect 288256 299950 288308 299956
rect 288164 248124 288216 248130
rect 288164 248066 288216 248072
rect 288072 248056 288124 248062
rect 288072 247998 288124 248004
rect 287888 247716 287940 247722
rect 287888 247658 287940 247664
rect 287900 247081 287928 247658
rect 288084 247081 288112 247998
rect 287886 247072 287942 247081
rect 287886 247007 287942 247016
rect 288070 247072 288126 247081
rect 288070 247007 288126 247016
rect 287612 159588 287664 159594
rect 287612 159530 287664 159536
rect 288176 158982 288204 248066
rect 288164 158976 288216 158982
rect 288164 158918 288216 158924
rect 288268 158506 288296 299950
rect 288348 244520 288400 244526
rect 288348 244462 288400 244468
rect 288256 158500 288308 158506
rect 288256 158442 288308 158448
rect 288268 157962 288296 158442
rect 288256 157956 288308 157962
rect 288256 157898 288308 157904
rect 287520 156596 287572 156602
rect 287520 156538 287572 156544
rect 287428 153876 287480 153882
rect 287428 153818 287480 153824
rect 287336 147008 287388 147014
rect 287336 146950 287388 146956
rect 287244 145716 287296 145722
rect 287244 145658 287296 145664
rect 287244 145580 287296 145586
rect 287244 145522 287296 145528
rect 287256 16574 287284 145522
rect 287256 16546 287376 16574
rect 287152 14476 287204 14482
rect 287152 14418 287204 14424
rect 287060 11756 287112 11762
rect 287060 11698 287112 11704
rect 286324 4888 286376 4894
rect 286324 4830 286376 4836
rect 286244 3454 286640 3482
rect 286612 480 286640 3454
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 288360 4146 288388 244462
rect 288452 131782 288480 306342
rect 288544 134570 288572 306410
rect 288636 305980 288664 310406
rect 288820 306474 288848 310420
rect 288808 306468 288860 306474
rect 288808 306410 288860 306416
rect 288636 305952 288756 305980
rect 288624 305584 288676 305590
rect 288624 305526 288676 305532
rect 288636 142934 288664 305526
rect 288728 144294 288756 305952
rect 288808 305516 288860 305522
rect 288808 305458 288860 305464
rect 288820 152658 288848 305458
rect 289004 292574 289032 310420
rect 289084 307828 289136 307834
rect 289084 307770 289136 307776
rect 288912 292546 289032 292574
rect 288912 155310 288940 292546
rect 288992 247512 289044 247518
rect 288992 247454 289044 247460
rect 289004 247081 289032 247454
rect 288990 247072 289046 247081
rect 288990 247007 289046 247016
rect 288900 155304 288952 155310
rect 288900 155246 288952 155252
rect 288808 152652 288860 152658
rect 288808 152594 288860 152600
rect 288716 144288 288768 144294
rect 288716 144230 288768 144236
rect 288624 142928 288676 142934
rect 288624 142870 288676 142876
rect 288532 134564 288584 134570
rect 288532 134506 288584 134512
rect 288440 131776 288492 131782
rect 288440 131718 288492 131724
rect 288992 6928 289044 6934
rect 288992 6870 289044 6876
rect 288348 4140 288400 4146
rect 288348 4082 288400 4088
rect 289004 480 289032 6870
rect 289096 6866 289124 307770
rect 289188 305590 289216 310420
rect 289280 310406 289478 310434
rect 289280 306406 289308 310406
rect 289268 306400 289320 306406
rect 289268 306342 289320 306348
rect 289176 305584 289228 305590
rect 289176 305526 289228 305532
rect 289648 305522 289676 310420
rect 289832 306406 289860 310420
rect 290016 310406 290122 310434
rect 289820 306400 289872 306406
rect 289820 306342 289872 306348
rect 290016 305674 290044 310406
rect 290292 309058 290320 310420
rect 290280 309052 290332 309058
rect 290280 308994 290332 309000
rect 290096 306400 290148 306406
rect 290096 306342 290148 306348
rect 289924 305646 290044 305674
rect 289636 305516 289688 305522
rect 289636 305458 289688 305464
rect 289820 305516 289872 305522
rect 289820 305458 289872 305464
rect 289544 305448 289596 305454
rect 289544 305390 289596 305396
rect 289176 247988 289228 247994
rect 289176 247930 289228 247936
rect 289188 247081 289216 247930
rect 289174 247072 289230 247081
rect 289174 247007 289230 247016
rect 289266 158808 289322 158817
rect 289266 158743 289322 158752
rect 289084 6860 289136 6866
rect 289084 6802 289136 6808
rect 289280 6594 289308 158743
rect 289450 155816 289506 155825
rect 289450 155751 289506 155760
rect 289358 153096 289414 153105
rect 289358 153031 289414 153040
rect 289268 6588 289320 6594
rect 289268 6530 289320 6536
rect 289372 6390 289400 153031
rect 289464 6458 289492 155751
rect 289556 155446 289584 305390
rect 289636 246696 289688 246702
rect 289636 246638 289688 246644
rect 289648 158914 289676 246638
rect 289728 244928 289780 244934
rect 289728 244870 289780 244876
rect 289636 158908 289688 158914
rect 289636 158850 289688 158856
rect 289634 155952 289690 155961
rect 289634 155887 289690 155896
rect 289544 155440 289596 155446
rect 289544 155382 289596 155388
rect 289556 154902 289584 155382
rect 289544 154896 289596 154902
rect 289544 154838 289596 154844
rect 289648 6526 289676 155887
rect 289636 6520 289688 6526
rect 289636 6462 289688 6468
rect 289452 6452 289504 6458
rect 289452 6394 289504 6400
rect 289360 6384 289412 6390
rect 289360 6326 289412 6332
rect 289740 3738 289768 244870
rect 289832 15910 289860 305458
rect 289924 130422 289952 305646
rect 290004 305584 290056 305590
rect 290004 305526 290056 305532
rect 290016 146946 290044 305526
rect 290108 151162 290136 306342
rect 290476 305590 290504 310420
rect 290568 310406 290766 310434
rect 290464 305584 290516 305590
rect 290464 305526 290516 305532
rect 290568 305522 290596 310406
rect 290556 305516 290608 305522
rect 290556 305458 290608 305464
rect 290936 303226 290964 310420
rect 291016 307964 291068 307970
rect 291016 307906 291068 307912
rect 290844 303198 290964 303226
rect 290844 302234 290872 303198
rect 290200 302206 290872 302234
rect 290200 156670 290228 302206
rect 290832 300688 290884 300694
rect 290832 300630 290884 300636
rect 290740 299940 290792 299946
rect 290740 299882 290792 299888
rect 290648 247920 290700 247926
rect 290648 247862 290700 247868
rect 290660 247081 290688 247862
rect 290646 247072 290702 247081
rect 290646 247007 290702 247016
rect 290752 158574 290780 299882
rect 290740 158568 290792 158574
rect 290740 158510 290792 158516
rect 290648 158500 290700 158506
rect 290648 158442 290700 158448
rect 290660 156806 290688 158442
rect 290752 157894 290780 158510
rect 290740 157888 290792 157894
rect 290740 157830 290792 157836
rect 290648 156800 290700 156806
rect 290648 156742 290700 156748
rect 290188 156664 290240 156670
rect 290188 156606 290240 156612
rect 290660 156330 290688 156742
rect 290738 156632 290794 156641
rect 290738 156567 290794 156576
rect 290648 156324 290700 156330
rect 290648 156266 290700 156272
rect 290096 151156 290148 151162
rect 290096 151098 290148 151104
rect 290004 146940 290056 146946
rect 290004 146882 290056 146888
rect 289912 130416 289964 130422
rect 289912 130358 289964 130364
rect 289820 15904 289872 15910
rect 289820 15846 289872 15852
rect 290752 6254 290780 156567
rect 290844 154426 290872 300630
rect 291028 292574 291056 307906
rect 291212 306406 291240 310420
rect 291200 306400 291252 306406
rect 291200 306342 291252 306348
rect 291200 305584 291252 305590
rect 291200 305526 291252 305532
rect 290936 292546 291056 292574
rect 290936 158506 290964 292546
rect 291016 245608 291068 245614
rect 291016 245550 291068 245556
rect 291028 245177 291056 245550
rect 291014 245168 291070 245177
rect 291014 245103 291070 245112
rect 291108 245064 291160 245070
rect 291108 245006 291160 245012
rect 291016 244996 291068 245002
rect 291016 244938 291068 244944
rect 290924 158500 290976 158506
rect 290924 158442 290976 158448
rect 290922 157992 290978 158001
rect 290922 157927 290978 157936
rect 290936 157282 290964 157927
rect 290924 157276 290976 157282
rect 290924 157218 290976 157224
rect 290922 156768 290978 156777
rect 290922 156703 290978 156712
rect 290832 154420 290884 154426
rect 290832 154362 290884 154368
rect 290936 6322 290964 156703
rect 291028 6662 291056 244938
rect 291016 6656 291068 6662
rect 291016 6598 291068 6604
rect 290924 6316 290976 6322
rect 290924 6258 290976 6264
rect 290740 6248 290792 6254
rect 290740 6190 290792 6196
rect 290188 4956 290240 4962
rect 290188 4898 290240 4904
rect 289728 3732 289780 3738
rect 289728 3674 289780 3680
rect 290200 480 290228 4898
rect 291120 3874 291148 245006
rect 291212 127634 291240 305526
rect 291396 304314 291424 310420
rect 291304 304286 291424 304314
rect 291304 129062 291332 304286
rect 291384 304224 291436 304230
rect 291384 304166 291436 304172
rect 291396 140078 291424 304166
rect 291488 141438 291516 310490
rect 291594 310406 291792 310434
rect 291568 306400 291620 306406
rect 291568 306342 291620 306348
rect 291660 306400 291712 306406
rect 291660 306342 291712 306348
rect 291580 148442 291608 306342
rect 291672 155242 291700 306342
rect 291764 244526 291792 310406
rect 292040 305590 292068 310420
rect 292224 306406 292252 310420
rect 292316 310406 292514 310434
rect 292212 306400 292264 306406
rect 292212 306342 292264 306348
rect 292028 305584 292080 305590
rect 292028 305526 292080 305532
rect 292316 304230 292344 310406
rect 292684 307834 292712 310420
rect 292672 307828 292724 307834
rect 292672 307770 292724 307776
rect 292672 306536 292724 306542
rect 292672 306478 292724 306484
rect 292580 306468 292632 306474
rect 292580 306410 292632 306416
rect 292304 304224 292356 304230
rect 292304 304166 292356 304172
rect 292304 300280 292356 300286
rect 292304 300222 292356 300228
rect 292212 245540 292264 245546
rect 292212 245482 292264 245488
rect 291752 244520 291804 244526
rect 291752 244462 291804 244468
rect 291752 244384 291804 244390
rect 291750 244352 291752 244361
rect 292224 244361 292252 245482
rect 291804 244352 291806 244361
rect 291750 244287 291806 244296
rect 292210 244352 292266 244361
rect 292210 244287 292266 244296
rect 292212 198076 292264 198082
rect 292212 198018 292264 198024
rect 292118 196072 292174 196081
rect 292118 196007 292174 196016
rect 291660 155236 291712 155242
rect 291660 155178 291712 155184
rect 291568 148436 291620 148442
rect 291568 148378 291620 148384
rect 291476 141432 291528 141438
rect 291476 141374 291528 141380
rect 291476 140208 291528 140214
rect 291476 140150 291528 140156
rect 291384 140072 291436 140078
rect 291384 140014 291436 140020
rect 291292 129056 291344 129062
rect 291292 128998 291344 129004
rect 291200 127628 291252 127634
rect 291200 127570 291252 127576
rect 291488 6914 291516 140150
rect 291396 6886 291516 6914
rect 291108 3868 291160 3874
rect 291108 3810 291160 3816
rect 291396 480 291424 6886
rect 292132 3398 292160 196007
rect 292224 158846 292252 198018
rect 292316 167006 292344 300222
rect 292488 248328 292540 248334
rect 292488 248270 292540 248276
rect 292396 247852 292448 247858
rect 292396 247794 292448 247800
rect 292408 247081 292436 247794
rect 292394 247072 292450 247081
rect 292394 247007 292450 247016
rect 292500 245290 292528 248270
rect 292408 245262 292528 245290
rect 292408 197334 292436 245262
rect 292488 245132 292540 245138
rect 292488 245074 292540 245080
rect 292396 197328 292448 197334
rect 292396 197270 292448 197276
rect 292304 167000 292356 167006
rect 292304 166942 292356 166948
rect 292394 166288 292450 166297
rect 292394 166223 292450 166232
rect 292212 158840 292264 158846
rect 292212 158782 292264 158788
rect 292408 6186 292436 166223
rect 292500 6730 292528 245074
rect 292592 17270 292620 306410
rect 292684 138718 292712 306478
rect 292776 145654 292804 310490
rect 292882 310406 293080 310434
rect 292856 306400 292908 306406
rect 292856 306342 292908 306348
rect 292868 149802 292896 306342
rect 293052 302234 293080 310406
rect 293224 308100 293276 308106
rect 293224 308042 293276 308048
rect 293052 302206 293172 302234
rect 293144 296714 293172 302206
rect 292960 296686 293172 296714
rect 292960 151094 292988 296686
rect 292948 151088 293000 151094
rect 292948 151030 293000 151036
rect 292856 149796 292908 149802
rect 292856 149738 292908 149744
rect 292764 145648 292816 145654
rect 292764 145590 292816 145596
rect 292672 138712 292724 138718
rect 292672 138654 292724 138660
rect 292580 17264 292632 17270
rect 292580 17206 292632 17212
rect 293236 16574 293264 308042
rect 293328 306474 293356 310420
rect 293420 310406 293618 310434
rect 293316 306468 293368 306474
rect 293316 306410 293368 306416
rect 293420 306406 293448 310406
rect 293500 309052 293552 309058
rect 293500 308994 293552 309000
rect 293408 306400 293460 306406
rect 293408 306342 293460 306348
rect 293512 302234 293540 308994
rect 293788 306542 293816 310420
rect 293972 307902 294000 310420
rect 293960 307896 294012 307902
rect 293960 307838 294012 307844
rect 293776 306536 293828 306542
rect 293776 306478 293828 306484
rect 294052 306536 294104 306542
rect 294052 306478 294104 306484
rect 293960 306468 294012 306474
rect 293960 306410 294012 306416
rect 293776 302864 293828 302870
rect 293776 302806 293828 302812
rect 293592 302728 293644 302734
rect 293592 302670 293644 302676
rect 293328 302206 293540 302234
rect 293328 159526 293356 302206
rect 293408 245404 293460 245410
rect 293408 245346 293460 245352
rect 293420 244497 293448 245346
rect 293406 244488 293462 244497
rect 293406 244423 293462 244432
rect 293316 159520 293368 159526
rect 293316 159462 293368 159468
rect 293498 158808 293554 158817
rect 293498 158743 293554 158752
rect 293236 16546 293356 16574
rect 293224 11824 293276 11830
rect 293224 11766 293276 11772
rect 292488 6724 292540 6730
rect 292488 6666 292540 6672
rect 292396 6180 292448 6186
rect 292396 6122 292448 6128
rect 292580 3528 292632 3534
rect 292580 3470 292632 3476
rect 292120 3392 292172 3398
rect 292120 3334 292172 3340
rect 292592 480 292620 3470
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 11766
rect 293328 3194 293356 16546
rect 293512 3670 293540 158743
rect 293604 158506 293632 302670
rect 293684 245472 293736 245478
rect 293684 245414 293736 245420
rect 293696 244361 293724 245414
rect 293682 244352 293738 244361
rect 293682 244287 293738 244296
rect 293684 243772 293736 243778
rect 293684 243714 293736 243720
rect 293696 159322 293724 243714
rect 293684 159316 293736 159322
rect 293684 159258 293736 159264
rect 293788 158710 293816 302806
rect 293866 158944 293922 158953
rect 293866 158879 293922 158888
rect 293776 158704 293828 158710
rect 293776 158646 293828 158652
rect 293592 158500 293644 158506
rect 293592 158442 293644 158448
rect 293500 3664 293552 3670
rect 293500 3606 293552 3612
rect 293880 3602 293908 158879
rect 293972 137290 294000 306410
rect 294064 144226 294092 306478
rect 294144 306400 294196 306406
rect 294144 306342 294196 306348
rect 294248 306354 294276 310420
rect 294432 306474 294460 310420
rect 294512 307828 294564 307834
rect 294512 307770 294564 307776
rect 294420 306468 294472 306474
rect 294420 306410 294472 306416
rect 294156 145586 294184 306342
rect 294248 306326 294368 306354
rect 294236 305516 294288 305522
rect 294236 305458 294288 305464
rect 294248 148374 294276 305458
rect 294340 152590 294368 306326
rect 294524 302234 294552 307770
rect 294616 306406 294644 310420
rect 294708 310406 294906 310434
rect 294604 306400 294656 306406
rect 294604 306342 294656 306348
rect 294708 305522 294736 310406
rect 295076 306542 295104 310420
rect 295260 307834 295288 310420
rect 295352 310406 295550 310434
rect 295734 310406 295932 310434
rect 295248 307828 295300 307834
rect 295248 307770 295300 307776
rect 295064 306536 295116 306542
rect 295064 306478 295116 306484
rect 294696 305516 294748 305522
rect 294696 305458 294748 305464
rect 295064 305312 295116 305318
rect 295064 305254 295116 305260
rect 294972 302796 295024 302802
rect 294972 302738 295024 302744
rect 294524 302206 294644 302234
rect 294328 152584 294380 152590
rect 294328 152526 294380 152532
rect 294236 148368 294288 148374
rect 294236 148310 294288 148316
rect 294144 145580 294196 145586
rect 294144 145522 294196 145528
rect 294052 144220 294104 144226
rect 294052 144162 294104 144168
rect 293960 137284 294012 137290
rect 293960 137226 294012 137232
rect 294616 126274 294644 302206
rect 294984 158574 295012 302738
rect 294972 158568 295024 158574
rect 294972 158510 295024 158516
rect 295076 158370 295104 305254
rect 295248 245336 295300 245342
rect 295248 245278 295300 245284
rect 295156 245200 295208 245206
rect 295156 245142 295208 245148
rect 295064 158364 295116 158370
rect 295064 158306 295116 158312
rect 295062 157448 295118 157457
rect 295062 157383 295118 157392
rect 294604 126268 294656 126274
rect 294604 126210 294656 126216
rect 294880 6792 294932 6798
rect 294880 6734 294932 6740
rect 293868 3596 293920 3602
rect 293868 3538 293920 3544
rect 293316 3188 293368 3194
rect 293316 3130 293368 3136
rect 294892 480 294920 6734
rect 295076 3534 295104 157383
rect 295168 3806 295196 245142
rect 295260 244769 295288 245278
rect 295246 244760 295302 244769
rect 295246 244695 295302 244704
rect 295248 244656 295300 244662
rect 295248 244598 295300 244604
rect 295260 3942 295288 244598
rect 295352 4078 295380 310406
rect 295800 307896 295852 307902
rect 295800 307838 295852 307844
rect 295432 306536 295484 306542
rect 295432 306478 295484 306484
rect 295340 4072 295392 4078
rect 295340 4014 295392 4020
rect 295444 4010 295472 306478
rect 295616 306468 295668 306474
rect 295616 306410 295668 306416
rect 295524 306400 295576 306406
rect 295524 306342 295576 306348
rect 295536 6798 295564 306342
rect 295628 142866 295656 306410
rect 295812 305522 295840 307838
rect 295800 305516 295852 305522
rect 295800 305458 295852 305464
rect 295904 296714 295932 310406
rect 295996 306406 296024 310420
rect 296076 307828 296128 307834
rect 296076 307770 296128 307776
rect 295984 306400 296036 306406
rect 295984 306342 296036 306348
rect 295984 305516 296036 305522
rect 295984 305458 296036 305464
rect 295720 296686 295932 296714
rect 295720 149734 295748 296686
rect 295708 149728 295760 149734
rect 295708 149670 295760 149676
rect 295616 142860 295668 142866
rect 295616 142802 295668 142808
rect 295996 29646 296024 305458
rect 296088 124914 296116 307770
rect 296180 306542 296208 310420
rect 296260 309052 296312 309058
rect 296260 308994 296312 309000
rect 296168 306536 296220 306542
rect 296168 306478 296220 306484
rect 296272 296714 296300 308994
rect 296364 306474 296392 310420
rect 296640 307873 296668 310420
rect 296626 307864 296682 307873
rect 296626 307799 296682 307808
rect 296352 306468 296404 306474
rect 296352 306410 296404 306416
rect 296720 306400 296772 306406
rect 296720 306342 296772 306348
rect 296628 300552 296680 300558
rect 296628 300494 296680 300500
rect 296180 296686 296300 296714
rect 296180 158778 296208 296686
rect 296536 246764 296588 246770
rect 296536 246706 296588 246712
rect 296548 159050 296576 246706
rect 296640 195974 296668 300494
rect 296732 244905 296760 306342
rect 296824 246265 296852 310420
rect 297008 308281 297036 310420
rect 296994 308272 297050 308281
rect 296994 308207 297050 308216
rect 297284 308009 297312 310420
rect 297270 308000 297326 308009
rect 297270 307935 297326 307944
rect 297468 306406 297496 310420
rect 297652 307873 297680 310420
rect 297928 308145 297956 310420
rect 298112 309097 298140 310420
rect 298204 310406 298402 310434
rect 298098 309088 298154 309097
rect 298098 309023 298154 309032
rect 297914 308136 297970 308145
rect 297914 308071 297970 308080
rect 297638 307864 297694 307873
rect 297638 307799 297694 307808
rect 297456 306400 297508 306406
rect 297456 306342 297508 306348
rect 298100 306400 298152 306406
rect 298100 306342 298152 306348
rect 298008 305244 298060 305250
rect 298008 305186 298060 305192
rect 297732 253360 297784 253366
rect 297732 253302 297784 253308
rect 297272 252068 297324 252074
rect 297272 252010 297324 252016
rect 297088 247580 297140 247586
rect 297088 247522 297140 247528
rect 296810 246256 296866 246265
rect 296810 246191 296866 246200
rect 296718 244896 296774 244905
rect 296718 244831 296774 244840
rect 296628 195968 296680 195974
rect 296628 195910 296680 195916
rect 297100 189961 297128 247522
rect 297180 246832 297232 246838
rect 297180 246774 297232 246780
rect 297192 198082 297220 246774
rect 297284 243574 297312 252010
rect 297364 247036 297416 247042
rect 297364 246978 297416 246984
rect 297272 243568 297324 243574
rect 297272 243510 297324 243516
rect 297180 198076 297232 198082
rect 297180 198018 297232 198024
rect 297284 195945 297312 243510
rect 297270 195936 297326 195945
rect 297270 195871 297326 195880
rect 297376 192817 297404 246978
rect 297456 246288 297508 246294
rect 297456 246230 297508 246236
rect 297362 192808 297418 192817
rect 297362 192743 297418 192752
rect 297270 191720 297326 191729
rect 297270 191655 297326 191664
rect 297284 191049 297312 191655
rect 297270 191040 297326 191049
rect 297270 190975 297326 190984
rect 297086 189952 297142 189961
rect 297086 189887 297142 189896
rect 297100 189145 297128 189887
rect 297086 189136 297142 189145
rect 297086 189071 297142 189080
rect 297180 171080 297232 171086
rect 297180 171022 297232 171028
rect 297192 169969 297220 171022
rect 297178 169960 297234 169969
rect 297178 169895 297234 169904
rect 296720 167000 296772 167006
rect 296720 166942 296772 166948
rect 296536 159044 296588 159050
rect 296536 158986 296588 158992
rect 296168 158772 296220 158778
rect 296168 158714 296220 158720
rect 296732 153610 296760 166942
rect 297284 159866 297312 190975
rect 297272 159860 297324 159866
rect 297272 159802 297324 159808
rect 297376 159798 297404 192743
rect 297468 191729 297496 246230
rect 297640 244724 297692 244730
rect 297640 244666 297692 244672
rect 297548 197464 297600 197470
rect 297548 197406 297600 197412
rect 297454 191720 297510 191729
rect 297454 191655 297510 191664
rect 297454 189136 297510 189145
rect 297454 189071 297510 189080
rect 297364 159792 297416 159798
rect 297364 159734 297416 159740
rect 297468 157690 297496 189071
rect 297560 159254 297588 197406
rect 297652 168065 297680 244666
rect 297744 168337 297772 253302
rect 297824 248260 297876 248266
rect 297824 248202 297876 248208
rect 297730 168328 297786 168337
rect 297730 168263 297786 168272
rect 297638 168056 297694 168065
rect 297638 167991 297694 168000
rect 297744 167686 297772 168263
rect 297732 167680 297784 167686
rect 297732 167622 297784 167628
rect 297548 159248 297600 159254
rect 297548 159190 297600 159196
rect 297836 158778 297864 248202
rect 297916 243568 297968 243574
rect 297916 243510 297968 243516
rect 297824 158772 297876 158778
rect 297824 158714 297876 158720
rect 297456 157684 297508 157690
rect 297456 157626 297508 157632
rect 297928 154494 297956 243510
rect 298020 158642 298048 305186
rect 298008 158636 298060 158642
rect 298008 158578 298060 158584
rect 298020 158234 298048 158578
rect 298008 158228 298060 158234
rect 298008 158170 298060 158176
rect 297916 154488 297968 154494
rect 297916 154430 297968 154436
rect 297456 154080 297508 154086
rect 297456 154022 297508 154028
rect 297468 153610 297496 154022
rect 296720 153604 296772 153610
rect 296720 153546 296772 153552
rect 297456 153604 297508 153610
rect 297456 153546 297508 153552
rect 296076 124908 296128 124914
rect 296076 124850 296128 124856
rect 295984 29640 296036 29646
rect 295984 29582 296036 29588
rect 298112 7614 298140 306342
rect 298204 159458 298232 310406
rect 298572 306406 298600 310420
rect 298560 306400 298612 306406
rect 298560 306342 298612 306348
rect 298756 302234 298784 310420
rect 299032 307873 299060 310420
rect 299216 308009 299244 310420
rect 299202 308000 299258 308009
rect 299202 307935 299258 307944
rect 299018 307864 299074 307873
rect 299018 307799 299074 307808
rect 298296 302206 298784 302234
rect 298192 159452 298244 159458
rect 298192 159394 298244 159400
rect 298296 159361 298324 302206
rect 299400 296714 299428 310420
rect 299572 306536 299624 306542
rect 299572 306478 299624 306484
rect 299480 306468 299532 306474
rect 299480 306410 299532 306416
rect 298388 296686 299428 296714
rect 298388 244361 298416 296686
rect 298836 248396 298888 248402
rect 298836 248338 298888 248344
rect 298744 247104 298796 247110
rect 298744 247046 298796 247052
rect 298756 244361 298784 247046
rect 298374 244352 298430 244361
rect 298374 244287 298430 244296
rect 298742 244352 298798 244361
rect 298742 244287 298798 244296
rect 298744 243500 298796 243506
rect 298744 243442 298796 243448
rect 298376 195968 298428 195974
rect 298376 195910 298428 195916
rect 298282 159352 298338 159361
rect 298282 159287 298338 159296
rect 298388 154970 298416 195910
rect 298756 188193 298784 243442
rect 298848 197470 298876 248338
rect 298928 246968 298980 246974
rect 298928 246910 298980 246916
rect 298940 243438 298968 246910
rect 299388 246900 299440 246906
rect 299388 246842 299440 246848
rect 299294 245576 299350 245585
rect 299294 245511 299350 245520
rect 299112 244860 299164 244866
rect 299112 244802 299164 244808
rect 299020 244792 299072 244798
rect 299020 244734 299072 244740
rect 299032 243506 299060 244734
rect 299020 243500 299072 243506
rect 299020 243442 299072 243448
rect 298928 243432 298980 243438
rect 298928 243374 298980 243380
rect 298836 197464 298888 197470
rect 298836 197406 298888 197412
rect 298836 197328 298888 197334
rect 298836 197270 298888 197276
rect 298742 188184 298798 188193
rect 298742 188119 298798 188128
rect 298848 159390 298876 197270
rect 298940 196897 298968 243374
rect 298926 196888 298982 196897
rect 298926 196823 298982 196832
rect 299124 193769 299152 244802
rect 299308 244390 299336 245511
rect 299296 244384 299348 244390
rect 299296 244326 299348 244332
rect 299296 243704 299348 243710
rect 299296 243646 299348 243652
rect 299204 243636 299256 243642
rect 299204 243578 299256 243584
rect 299110 193760 299166 193769
rect 299110 193695 299166 193704
rect 299124 190454 299152 193695
rect 298940 190426 299152 190454
rect 298940 159934 298968 190426
rect 299110 187776 299166 187785
rect 299110 187711 299166 187720
rect 298928 159928 298980 159934
rect 298928 159870 298980 159876
rect 298836 159384 298888 159390
rect 298836 159326 298888 159332
rect 299018 158808 299074 158817
rect 299018 158743 299074 158752
rect 298376 154964 298428 154970
rect 298376 154906 298428 154912
rect 299032 8974 299060 158743
rect 299124 152522 299152 187711
rect 299216 158302 299244 243578
rect 299308 158930 299336 243646
rect 299400 159118 299428 246842
rect 299492 244662 299520 306410
rect 299584 245138 299612 306478
rect 299572 245132 299624 245138
rect 299572 245074 299624 245080
rect 299676 245070 299704 310420
rect 299756 306400 299808 306406
rect 299756 306342 299808 306348
rect 299860 306354 299888 310420
rect 300044 306474 300072 310420
rect 300136 310406 300334 310434
rect 300136 306542 300164 310406
rect 300124 306536 300176 306542
rect 300124 306478 300176 306484
rect 300032 306468 300084 306474
rect 300032 306410 300084 306416
rect 299664 245064 299716 245070
rect 299664 245006 299716 245012
rect 299480 244656 299532 244662
rect 299768 244633 299796 306342
rect 299860 306326 299980 306354
rect 299848 305516 299900 305522
rect 299848 305458 299900 305464
rect 299860 248169 299888 305458
rect 299846 248160 299902 248169
rect 299846 248095 299902 248104
rect 299952 248033 299980 306326
rect 300504 305522 300532 310420
rect 300596 310406 300794 310434
rect 300596 306406 300624 310406
rect 300584 306400 300636 306406
rect 300584 306342 300636 306348
rect 300492 305516 300544 305522
rect 300492 305458 300544 305464
rect 299938 248024 299994 248033
rect 299938 247959 299994 247968
rect 300674 248024 300730 248033
rect 300674 247959 300730 247968
rect 300688 247722 300716 247959
rect 300676 247716 300728 247722
rect 300676 247658 300728 247664
rect 300768 247648 300820 247654
rect 300768 247590 300820 247596
rect 299480 244598 299532 244604
rect 299754 244624 299810 244633
rect 299754 244559 299810 244568
rect 300780 243778 300808 247590
rect 300872 245206 300900 310490
rect 300964 306354 300992 310420
rect 301162 310406 301360 310434
rect 301228 306400 301280 306406
rect 300964 306326 301176 306354
rect 301228 306342 301280 306348
rect 300952 305516 301004 305522
rect 300952 305458 301004 305464
rect 300964 245313 300992 305458
rect 301044 305448 301096 305454
rect 301044 305390 301096 305396
rect 300950 245304 301006 245313
rect 300950 245239 301006 245248
rect 300860 245200 300912 245206
rect 300860 245142 300912 245148
rect 301056 244769 301084 305390
rect 301148 245002 301176 306326
rect 301240 247625 301268 306342
rect 301226 247616 301282 247625
rect 301226 247551 301282 247560
rect 301332 247353 301360 310406
rect 301608 305522 301636 310420
rect 301792 306406 301820 310420
rect 301884 310406 302082 310434
rect 301780 306400 301832 306406
rect 301780 306342 301832 306348
rect 301596 305516 301648 305522
rect 301596 305458 301648 305464
rect 301884 305454 301912 310406
rect 302252 308360 302280 310420
rect 302450 310406 302648 310434
rect 302160 308332 302280 308360
rect 302160 307986 302188 308332
rect 302160 307958 302372 307986
rect 302240 306468 302292 306474
rect 302240 306410 302292 306416
rect 301872 305448 301924 305454
rect 301872 305390 301924 305396
rect 301318 247344 301374 247353
rect 301318 247279 301374 247288
rect 301136 244996 301188 245002
rect 301136 244938 301188 244944
rect 302252 244934 302280 306410
rect 302344 245449 302372 307958
rect 302424 306536 302476 306542
rect 302424 306478 302476 306484
rect 302330 245440 302386 245449
rect 302330 245375 302386 245384
rect 302436 245177 302464 306478
rect 302516 306400 302568 306406
rect 302516 306342 302568 306348
rect 302422 245168 302478 245177
rect 302422 245103 302478 245112
rect 302528 245041 302556 306342
rect 302620 247761 302648 310406
rect 302712 306474 302740 310420
rect 302700 306468 302752 306474
rect 302700 306410 302752 306416
rect 302896 306406 302924 310420
rect 302988 310406 303186 310434
rect 302884 306400 302936 306406
rect 302884 306342 302936 306348
rect 302988 302234 303016 310406
rect 303356 306542 303384 310420
rect 303344 306536 303396 306542
rect 303344 306478 303396 306484
rect 302712 302206 303016 302234
rect 302606 247752 302662 247761
rect 302606 247687 302662 247696
rect 302712 247489 302740 302206
rect 303540 296714 303568 310420
rect 303816 306610 303844 310420
rect 303804 306604 303856 306610
rect 303804 306546 303856 306552
rect 304000 306490 304028 310420
rect 302804 296686 303568 296714
rect 303632 306462 304028 306490
rect 302804 247897 302832 296686
rect 302790 247888 302846 247897
rect 302790 247823 302846 247832
rect 302698 247480 302754 247489
rect 302698 247415 302754 247424
rect 303632 245410 303660 306462
rect 303712 306400 303764 306406
rect 304184 306354 304212 310420
rect 303712 306342 303764 306348
rect 303724 245478 303752 306342
rect 303908 306326 304212 306354
rect 304276 310406 304474 310434
rect 303804 305380 303856 305386
rect 303804 305322 303856 305328
rect 303816 247518 303844 305322
rect 303908 247994 303936 306326
rect 304276 302234 304304 310406
rect 304356 306604 304408 306610
rect 304356 306546 304408 306552
rect 304000 302206 304304 302234
rect 303896 247988 303948 247994
rect 303896 247930 303948 247936
rect 303804 247512 303856 247518
rect 303804 247454 303856 247460
rect 304000 247450 304028 302206
rect 304368 296714 304396 306546
rect 304644 306406 304672 310420
rect 304632 306400 304684 306406
rect 304632 306342 304684 306348
rect 304828 305386 304856 310420
rect 305104 309134 305132 310420
rect 304920 309106 305132 309134
rect 304816 305380 304868 305386
rect 304816 305322 304868 305328
rect 304920 304298 304948 309106
rect 305288 306626 305316 310420
rect 305012 306598 305316 306626
rect 305380 310406 305578 310434
rect 304908 304292 304960 304298
rect 304908 304234 304960 304240
rect 304092 296686 304396 296714
rect 303988 247444 304040 247450
rect 303988 247386 304040 247392
rect 304092 247110 304120 296686
rect 304080 247104 304132 247110
rect 304080 247046 304132 247052
rect 303712 245472 303764 245478
rect 303712 245414 303764 245420
rect 303620 245404 303672 245410
rect 303620 245346 303672 245352
rect 305012 245342 305040 306598
rect 305380 306490 305408 310406
rect 305748 309134 305776 310420
rect 305196 306462 305408 306490
rect 305472 309106 305776 309134
rect 305092 305312 305144 305318
rect 305092 305254 305144 305260
rect 305104 245546 305132 305254
rect 305196 247926 305224 306462
rect 305276 305380 305328 305386
rect 305276 305322 305328 305328
rect 305288 248033 305316 305322
rect 305472 304450 305500 309106
rect 305932 305318 305960 310420
rect 306024 310406 306222 310434
rect 306024 305386 306052 310406
rect 306392 305386 306420 310420
rect 306590 310406 306696 310434
rect 306472 306468 306524 306474
rect 306472 306410 306524 306416
rect 306012 305380 306064 305386
rect 306012 305322 306064 305328
rect 306380 305380 306432 305386
rect 306380 305322 306432 305328
rect 305920 305312 305972 305318
rect 305920 305254 305972 305260
rect 306380 305244 306432 305250
rect 306380 305186 306432 305192
rect 305380 304422 305500 304450
rect 305274 248024 305330 248033
rect 305274 247959 305330 247968
rect 305184 247920 305236 247926
rect 305184 247862 305236 247868
rect 305380 247858 305408 304422
rect 305460 304292 305512 304298
rect 305460 304234 305512 304240
rect 305472 248062 305500 304234
rect 305460 248056 305512 248062
rect 305460 247998 305512 248004
rect 305368 247852 305420 247858
rect 305368 247794 305420 247800
rect 305092 245540 305144 245546
rect 305092 245482 305144 245488
rect 305000 245336 305052 245342
rect 305000 245278 305052 245284
rect 302514 245032 302570 245041
rect 302514 244967 302570 244976
rect 306392 244934 306420 305186
rect 306484 245206 306512 306410
rect 306564 306400 306616 306406
rect 306564 306342 306616 306348
rect 306576 245585 306604 306342
rect 306668 245614 306696 310406
rect 306760 310406 306866 310434
rect 306760 306474 306788 310406
rect 306748 306468 306800 306474
rect 306748 306410 306800 306416
rect 307036 306354 307064 310420
rect 307220 306406 307248 310420
rect 307312 310406 307510 310434
rect 306760 306326 307064 306354
rect 307208 306400 307260 306406
rect 307208 306342 307260 306348
rect 306656 245608 306708 245614
rect 306562 245576 306618 245585
rect 306656 245550 306708 245556
rect 306562 245511 306618 245520
rect 306472 245200 306524 245206
rect 306472 245142 306524 245148
rect 306760 245002 306788 306326
rect 306840 305380 306892 305386
rect 306840 305322 306892 305328
rect 306852 245274 306880 305322
rect 307312 305250 307340 310406
rect 307300 305244 307352 305250
rect 307300 305186 307352 305192
rect 307680 296714 307708 310420
rect 307864 310406 307970 310434
rect 307760 306400 307812 306406
rect 307760 306342 307812 306348
rect 306944 296686 307708 296714
rect 306944 248062 306972 296686
rect 306932 248056 306984 248062
rect 306932 247998 306984 248004
rect 306840 245268 306892 245274
rect 306840 245210 306892 245216
rect 307772 245070 307800 306342
rect 307864 245410 307892 310406
rect 308140 306354 308168 310420
rect 307956 306326 308168 306354
rect 307956 245546 307984 306326
rect 308036 305380 308088 305386
rect 308036 305322 308088 305328
rect 307944 245540 307996 245546
rect 307944 245482 307996 245488
rect 307852 245404 307904 245410
rect 307852 245346 307904 245352
rect 308048 245138 308076 305322
rect 308128 305312 308180 305318
rect 308128 305254 308180 305260
rect 308140 247625 308168 305254
rect 308324 296714 308352 310420
rect 308416 310406 308614 310434
rect 308416 306406 308444 310406
rect 308404 306400 308456 306406
rect 308404 306342 308456 306348
rect 308784 305386 308812 310420
rect 308772 305380 308824 305386
rect 308772 305322 308824 305328
rect 308968 305318 308996 310420
rect 309140 306400 309192 306406
rect 309140 306342 309192 306348
rect 308956 305312 309008 305318
rect 308956 305254 309008 305260
rect 308232 296686 308352 296714
rect 308232 247994 308260 296686
rect 308220 247988 308272 247994
rect 308220 247930 308272 247936
rect 308126 247616 308182 247625
rect 308126 247551 308182 247560
rect 309152 245342 309180 306342
rect 309244 306218 309272 310420
rect 309428 306490 309456 310420
rect 309428 306462 309548 306490
rect 309244 306190 309456 306218
rect 309324 305380 309376 305386
rect 309324 305322 309376 305328
rect 309232 305312 309284 305318
rect 309232 305254 309284 305260
rect 309140 245336 309192 245342
rect 309244 245313 309272 305254
rect 309336 245478 309364 305322
rect 309428 245614 309456 306190
rect 309520 305318 309548 306462
rect 309508 305312 309560 305318
rect 309508 305254 309560 305260
rect 309612 302234 309640 310420
rect 309704 310406 309902 310434
rect 309704 305386 309732 310406
rect 310072 306406 310100 310420
rect 310164 310406 310362 310434
rect 310060 306400 310112 306406
rect 310060 306342 310112 306348
rect 309692 305380 309744 305386
rect 309692 305322 309744 305328
rect 309520 302206 309640 302234
rect 309520 247926 309548 302206
rect 310164 296714 310192 310406
rect 310532 305386 310560 310420
rect 310520 305380 310572 305386
rect 310520 305322 310572 305328
rect 310520 305244 310572 305250
rect 310520 305186 310572 305192
rect 309612 296686 310192 296714
rect 309612 264450 309640 296686
rect 309600 264444 309652 264450
rect 309600 264386 309652 264392
rect 310532 250714 310560 305186
rect 310624 264382 310652 310490
rect 310730 310406 310836 310434
rect 310808 309134 310836 310406
rect 310808 309106 311020 309134
rect 310704 306400 310756 306406
rect 310704 306342 310756 306348
rect 310716 275466 310744 306342
rect 310888 305380 310940 305386
rect 310888 305322 310940 305328
rect 310796 304292 310848 304298
rect 310796 304234 310848 304240
rect 310808 276758 310836 304234
rect 310900 287745 310928 305322
rect 310992 298761 311020 309106
rect 311176 304298 311204 310420
rect 311360 305250 311388 310420
rect 311348 305244 311400 305250
rect 311348 305186 311400 305192
rect 311164 304292 311216 304298
rect 311164 304234 311216 304240
rect 311636 302977 311664 310420
rect 311820 306406 311848 310420
rect 311808 306400 311860 306406
rect 312004 306354 312032 310420
rect 312280 306474 312308 310420
rect 312268 306468 312320 306474
rect 312268 306410 312320 306416
rect 312464 306354 312492 310420
rect 311808 306342 311860 306348
rect 311912 306326 312032 306354
rect 312096 306326 312492 306354
rect 312556 310406 312754 310434
rect 311622 302968 311678 302977
rect 311622 302903 311678 302912
rect 310978 298752 311034 298761
rect 310978 298687 311034 298696
rect 310886 287736 310942 287745
rect 310886 287671 310942 287680
rect 310796 276752 310848 276758
rect 310796 276694 310848 276700
rect 310704 275460 310756 275466
rect 310704 275402 310756 275408
rect 310612 264376 310664 264382
rect 310612 264318 310664 264324
rect 310520 250708 310572 250714
rect 310520 250650 310572 250656
rect 311912 250646 311940 306326
rect 311992 305380 312044 305386
rect 311992 305322 312044 305328
rect 312004 271250 312032 305322
rect 312096 274174 312124 306326
rect 312556 306218 312584 310406
rect 312636 306468 312688 306474
rect 312636 306410 312688 306416
rect 312188 306190 312584 306218
rect 312188 287842 312216 306190
rect 312648 305969 312676 306410
rect 312634 305960 312690 305969
rect 312634 305895 312690 305904
rect 312924 302234 312952 310420
rect 313108 305386 313136 310420
rect 313280 306468 313332 306474
rect 313280 306410 313332 306416
rect 313096 305380 313148 305386
rect 313096 305322 313148 305328
rect 312280 302206 312952 302234
rect 312176 287836 312228 287842
rect 312176 287778 312228 287784
rect 312280 287774 312308 302206
rect 312268 287768 312320 287774
rect 312268 287710 312320 287716
rect 312084 274168 312136 274174
rect 312084 274110 312136 274116
rect 311992 271244 312044 271250
rect 311992 271186 312044 271192
rect 311900 250640 311952 250646
rect 311900 250582 311952 250588
rect 313292 249218 313320 306410
rect 313384 258806 313412 310420
rect 313464 306400 313516 306406
rect 313464 306342 313516 306348
rect 313476 269958 313504 306342
rect 313568 305538 313596 310420
rect 313752 306542 313780 310420
rect 313844 310406 314042 310434
rect 313740 306536 313792 306542
rect 313740 306478 313792 306484
rect 313568 305510 313780 305538
rect 313556 305380 313608 305386
rect 313556 305322 313608 305328
rect 313568 283762 313596 305322
rect 313648 304292 313700 304298
rect 313648 304234 313700 304240
rect 313660 284986 313688 304234
rect 313752 298994 313780 305510
rect 313844 305386 313872 310406
rect 313924 306536 313976 306542
rect 313924 306478 313976 306484
rect 313832 305380 313884 305386
rect 313832 305322 313884 305328
rect 313936 304298 313964 306478
rect 314212 306474 314240 310420
rect 314200 306468 314252 306474
rect 314200 306410 314252 306416
rect 314396 306406 314424 310420
rect 314672 306490 314700 310420
rect 314856 307834 314884 310420
rect 314844 307828 314896 307834
rect 314844 307770 314896 307776
rect 314672 306462 315068 306490
rect 314384 306400 314436 306406
rect 314384 306342 314436 306348
rect 314844 306400 314896 306406
rect 314844 306342 314896 306348
rect 314752 305312 314804 305318
rect 314752 305254 314804 305260
rect 314660 305244 314712 305250
rect 314660 305186 314712 305192
rect 313924 304292 313976 304298
rect 313924 304234 313976 304240
rect 313740 298988 313792 298994
rect 313740 298930 313792 298936
rect 313648 284980 313700 284986
rect 313648 284922 313700 284928
rect 313556 283756 313608 283762
rect 313556 283698 313608 283704
rect 313464 269952 313516 269958
rect 313464 269894 313516 269900
rect 313372 258800 313424 258806
rect 313372 258742 313424 258748
rect 313280 249212 313332 249218
rect 313280 249154 313332 249160
rect 314672 249150 314700 305186
rect 314764 263022 314792 305254
rect 314856 264314 314884 306342
rect 314936 305380 314988 305386
rect 314936 305322 314988 305328
rect 314948 268530 314976 305322
rect 315040 282266 315068 306462
rect 315132 302234 315160 310420
rect 315316 306406 315344 310420
rect 315304 306400 315356 306406
rect 315304 306342 315356 306348
rect 315500 305318 315528 310420
rect 315592 310406 315790 310434
rect 315592 305386 315620 310406
rect 315580 305380 315632 305386
rect 315580 305322 315632 305328
rect 315488 305312 315540 305318
rect 315488 305254 315540 305260
rect 315960 305250 315988 310420
rect 316144 307873 316172 310420
rect 316328 310406 316434 310434
rect 316130 307864 316186 307873
rect 316130 307799 316186 307808
rect 316132 306536 316184 306542
rect 316132 306478 316184 306484
rect 316040 306468 316092 306474
rect 316040 306410 316092 306416
rect 315948 305244 316000 305250
rect 315948 305186 316000 305192
rect 315132 302206 315436 302234
rect 315408 296714 315436 302206
rect 315132 296686 315436 296714
rect 315132 286550 315160 296686
rect 315120 286544 315172 286550
rect 315120 286486 315172 286492
rect 315028 282260 315080 282266
rect 315028 282202 315080 282208
rect 314936 268524 314988 268530
rect 314936 268466 314988 268472
rect 314844 264308 314896 264314
rect 314844 264250 314896 264256
rect 314752 263016 314804 263022
rect 314752 262958 314804 262964
rect 316052 254726 316080 306410
rect 316144 280906 316172 306478
rect 316224 306400 316276 306406
rect 316224 306342 316276 306348
rect 316236 294778 316264 306342
rect 316328 296070 316356 310406
rect 316604 304502 316632 310420
rect 316788 306474 316816 310420
rect 316880 310406 317078 310434
rect 316776 306468 316828 306474
rect 316776 306410 316828 306416
rect 316880 306406 316908 310406
rect 317248 306542 317276 310420
rect 317524 307902 317552 310420
rect 317512 307896 317564 307902
rect 317512 307838 317564 307844
rect 317236 306536 317288 306542
rect 317708 306490 317736 310420
rect 317236 306478 317288 306484
rect 317524 306462 317736 306490
rect 316868 306400 316920 306406
rect 316868 306342 316920 306348
rect 317420 306400 317472 306406
rect 317420 306342 317472 306348
rect 316592 304496 316644 304502
rect 316592 304438 316644 304444
rect 316316 296064 316368 296070
rect 316316 296006 316368 296012
rect 316224 294772 316276 294778
rect 316224 294714 316276 294720
rect 316132 280900 316184 280906
rect 316132 280842 316184 280848
rect 316040 254720 316092 254726
rect 316040 254662 316092 254668
rect 317432 254658 317460 306342
rect 317524 267102 317552 306462
rect 317892 306354 317920 310420
rect 317984 310406 318182 310434
rect 317984 306406 318012 310406
rect 318154 307864 318210 307873
rect 318064 307828 318116 307834
rect 318154 307799 318210 307808
rect 318064 307770 318116 307776
rect 317616 306326 317920 306354
rect 317972 306400 318024 306406
rect 317972 306342 318024 306348
rect 317616 278186 317644 306326
rect 317696 305380 317748 305386
rect 317696 305322 317748 305328
rect 317708 283694 317736 305322
rect 317696 283688 317748 283694
rect 317696 283630 317748 283636
rect 318076 282334 318104 307770
rect 318168 286482 318196 307799
rect 318352 307154 318380 310420
rect 318340 307148 318392 307154
rect 318340 307090 318392 307096
rect 318536 305386 318564 310420
rect 318812 305386 318840 310420
rect 318892 306400 318944 306406
rect 318996 306377 319024 310420
rect 318892 306342 318944 306348
rect 318982 306368 319038 306377
rect 318524 305380 318576 305386
rect 318524 305322 318576 305328
rect 318800 305380 318852 305386
rect 318800 305322 318852 305328
rect 318800 303748 318852 303754
rect 318800 303690 318852 303696
rect 318156 286476 318208 286482
rect 318156 286418 318208 286424
rect 318064 282328 318116 282334
rect 318064 282270 318116 282276
rect 317604 278180 317656 278186
rect 317604 278122 317656 278128
rect 317512 267096 317564 267102
rect 317512 267038 317564 267044
rect 318812 262954 318840 303690
rect 318904 265810 318932 306342
rect 318982 306303 319038 306312
rect 319180 305538 319208 310420
rect 319088 305510 319208 305538
rect 319272 310406 319470 310434
rect 318984 304292 319036 304298
rect 318984 304234 319036 304240
rect 318996 279546 319024 304234
rect 319088 282198 319116 305510
rect 319168 305380 319220 305386
rect 319168 305322 319220 305328
rect 319180 286414 319208 305322
rect 319272 304298 319300 310406
rect 319640 304434 319668 310420
rect 319824 306406 319852 310420
rect 319916 310406 320114 310434
rect 319812 306400 319864 306406
rect 319812 306342 319864 306348
rect 319628 304428 319680 304434
rect 319628 304370 319680 304376
rect 319260 304292 319312 304298
rect 319260 304234 319312 304240
rect 319916 303754 319944 310406
rect 320180 308236 320232 308242
rect 320180 308178 320232 308184
rect 320086 306368 320142 306377
rect 320086 306303 320142 306312
rect 320100 305833 320128 306303
rect 320086 305824 320142 305833
rect 320086 305759 320142 305768
rect 319904 303748 319956 303754
rect 319904 303690 319956 303696
rect 319168 286408 319220 286414
rect 319168 286350 319220 286356
rect 319076 282192 319128 282198
rect 319076 282134 319128 282140
rect 318984 279540 319036 279546
rect 318984 279482 319036 279488
rect 318892 265804 318944 265810
rect 318892 265746 318944 265752
rect 318800 262948 318852 262954
rect 318800 262890 318852 262896
rect 320192 261662 320220 308178
rect 320284 306678 320312 310420
rect 320376 310406 320574 310434
rect 320272 306672 320324 306678
rect 320272 306614 320324 306620
rect 320272 306536 320324 306542
rect 320272 306478 320324 306484
rect 320284 262886 320312 306478
rect 320376 264246 320404 310406
rect 320744 308242 320772 310420
rect 320732 308236 320784 308242
rect 320732 308178 320784 308184
rect 320928 308122 320956 310420
rect 320560 308094 320956 308122
rect 321020 310406 321218 310434
rect 320456 306400 320508 306406
rect 320456 306342 320508 306348
rect 320468 276690 320496 306342
rect 320560 301646 320588 308094
rect 320824 307896 320876 307902
rect 320824 307838 320876 307844
rect 320548 301640 320600 301646
rect 320548 301582 320600 301588
rect 320836 280974 320864 307838
rect 321020 306542 321048 310406
rect 321100 306672 321152 306678
rect 321100 306614 321152 306620
rect 321008 306536 321060 306542
rect 321008 306478 321060 306484
rect 321112 302841 321140 306614
rect 321388 306406 321416 310420
rect 321376 306400 321428 306406
rect 321376 306342 321428 306348
rect 321572 305386 321600 310420
rect 321664 310406 321862 310434
rect 321560 305380 321612 305386
rect 321560 305322 321612 305328
rect 321560 305244 321612 305250
rect 321560 305186 321612 305192
rect 321098 302832 321154 302841
rect 321098 302767 321154 302776
rect 320824 280968 320876 280974
rect 320824 280910 320876 280916
rect 320456 276684 320508 276690
rect 320456 276626 320508 276632
rect 320364 264240 320416 264246
rect 320364 264182 320416 264188
rect 320272 262880 320324 262886
rect 320272 262822 320324 262828
rect 320180 261656 320232 261662
rect 320180 261598 320232 261604
rect 317420 254652 317472 254658
rect 317420 254594 317472 254600
rect 321572 250578 321600 305186
rect 321664 261594 321692 310406
rect 322032 306354 322060 310420
rect 322216 307086 322244 310420
rect 322308 310406 322506 310434
rect 322204 307080 322256 307086
rect 322204 307022 322256 307028
rect 321756 306326 322060 306354
rect 321756 275398 321784 306326
rect 322308 306218 322336 310406
rect 321848 306190 322336 306218
rect 321848 280838 321876 306190
rect 321928 305380 321980 305386
rect 321928 305322 321980 305328
rect 321940 300121 321968 305322
rect 322676 305250 322704 310420
rect 322952 306474 322980 310420
rect 322940 306468 322992 306474
rect 322940 306410 322992 306416
rect 323136 306354 323164 310420
rect 323320 306490 323348 310420
rect 322952 306326 323164 306354
rect 323228 306462 323348 306490
rect 323412 310406 323610 310434
rect 322664 305244 322716 305250
rect 322664 305186 322716 305192
rect 321926 300112 321982 300121
rect 321926 300047 321982 300056
rect 321836 280832 321888 280838
rect 321836 280774 321888 280780
rect 321744 275392 321796 275398
rect 321744 275334 321796 275340
rect 321652 261588 321704 261594
rect 321652 261530 321704 261536
rect 321560 250572 321612 250578
rect 321560 250514 321612 250520
rect 314660 249144 314712 249150
rect 314660 249086 314712 249092
rect 309508 247920 309560 247926
rect 309508 247862 309560 247868
rect 322952 247858 322980 306326
rect 323228 306218 323256 306462
rect 323412 306354 323440 310406
rect 323492 306468 323544 306474
rect 323492 306410 323544 306416
rect 323136 306190 323256 306218
rect 323320 306326 323440 306354
rect 323032 305312 323084 305318
rect 323032 305254 323084 305260
rect 323044 252006 323072 305254
rect 323136 274106 323164 306190
rect 323216 305380 323268 305386
rect 323216 305322 323268 305328
rect 323228 278118 323256 305322
rect 323320 297566 323348 306326
rect 323504 302234 323532 306410
rect 323780 305386 323808 310420
rect 323768 305380 323820 305386
rect 323768 305322 323820 305328
rect 323964 305318 323992 310420
rect 324240 305697 324268 310420
rect 324320 306400 324372 306406
rect 324320 306342 324372 306348
rect 324226 305688 324282 305697
rect 324226 305623 324282 305632
rect 323952 305312 324004 305318
rect 323952 305254 324004 305260
rect 323412 302206 323532 302234
rect 323412 298926 323440 302206
rect 323400 298920 323452 298926
rect 323400 298862 323452 298868
rect 323308 297560 323360 297566
rect 323308 297502 323360 297508
rect 323216 278112 323268 278118
rect 323216 278054 323268 278060
rect 323124 274100 323176 274106
rect 323124 274042 323176 274048
rect 323032 252000 323084 252006
rect 323032 251942 323084 251948
rect 322940 247852 322992 247858
rect 322940 247794 322992 247800
rect 309416 245608 309468 245614
rect 309416 245550 309468 245556
rect 309324 245472 309376 245478
rect 309324 245414 309376 245420
rect 309140 245278 309192 245284
rect 309230 245304 309286 245313
rect 309230 245239 309286 245248
rect 324332 245177 324360 306342
rect 324424 305561 324452 310420
rect 324608 305674 324636 310420
rect 324516 305646 324636 305674
rect 324700 310406 324898 310434
rect 324410 305552 324466 305561
rect 324410 305487 324466 305496
rect 324412 305380 324464 305386
rect 324412 305322 324464 305328
rect 324424 247790 324452 305322
rect 324516 251938 324544 305646
rect 324594 305552 324650 305561
rect 324594 305487 324650 305496
rect 324608 279478 324636 305487
rect 324700 296002 324728 310406
rect 325068 306406 325096 310420
rect 325160 310406 325358 310434
rect 325056 306400 325108 306406
rect 325056 306342 325108 306348
rect 325160 305386 325188 310406
rect 325148 305380 325200 305386
rect 325148 305322 325200 305328
rect 325528 304366 325556 310420
rect 325726 310406 325924 310434
rect 325792 306604 325844 306610
rect 325792 306546 325844 306552
rect 325700 306468 325752 306474
rect 325700 306410 325752 306416
rect 325516 304360 325568 304366
rect 325516 304302 325568 304308
rect 324688 295996 324740 296002
rect 324688 295938 324740 295944
rect 324596 279472 324648 279478
rect 324596 279414 324648 279420
rect 324504 251932 324556 251938
rect 324504 251874 324556 251880
rect 324412 247784 324464 247790
rect 324412 247726 324464 247732
rect 324318 245168 324374 245177
rect 308036 245132 308088 245138
rect 324318 245103 324374 245112
rect 308036 245074 308088 245080
rect 307760 245064 307812 245070
rect 325712 245041 325740 306410
rect 325804 246566 325832 306546
rect 325896 306542 325924 310406
rect 325884 306536 325936 306542
rect 325884 306478 325936 306484
rect 325884 306400 325936 306406
rect 325884 306342 325936 306348
rect 325988 306354 326016 310420
rect 326172 306474 326200 310420
rect 326252 306536 326304 306542
rect 326252 306478 326304 306484
rect 326160 306468 326212 306474
rect 326160 306410 326212 306416
rect 325896 246634 325924 306342
rect 325988 306326 326200 306354
rect 325976 305380 326028 305386
rect 325976 305322 326028 305328
rect 325988 256018 326016 305322
rect 326068 305312 326120 305318
rect 326068 305254 326120 305260
rect 326080 257446 326108 305254
rect 326172 272610 326200 306326
rect 326264 298858 326292 306478
rect 326356 305386 326384 310420
rect 326448 310406 326646 310434
rect 326448 306406 326476 310406
rect 326816 306610 326844 310420
rect 326804 306604 326856 306610
rect 326804 306546 326856 306552
rect 326436 306400 326488 306406
rect 326436 306342 326488 306348
rect 326344 305380 326396 305386
rect 326344 305322 326396 305328
rect 327000 305318 327028 310420
rect 327172 306536 327224 306542
rect 327172 306478 327224 306484
rect 327080 306468 327132 306474
rect 327080 306410 327132 306416
rect 326988 305312 327040 305318
rect 326988 305254 327040 305260
rect 326252 298852 326304 298858
rect 326252 298794 326304 298800
rect 326160 272604 326212 272610
rect 326160 272546 326212 272552
rect 326068 257440 326120 257446
rect 326068 257382 326120 257388
rect 325976 256012 326028 256018
rect 325976 255954 326028 255960
rect 325884 246628 325936 246634
rect 325884 246570 325936 246576
rect 325792 246560 325844 246566
rect 325792 246502 325844 246508
rect 307760 245006 307812 245012
rect 325698 245032 325754 245041
rect 306748 244996 306800 245002
rect 325698 244967 325754 244976
rect 306748 244938 306800 244944
rect 302240 244928 302292 244934
rect 302240 244870 302292 244876
rect 306380 244928 306432 244934
rect 327092 244905 327120 306410
rect 327184 246498 327212 306478
rect 327276 269890 327304 310420
rect 327368 275330 327396 310490
rect 327474 310406 327672 310434
rect 327448 306400 327500 306406
rect 327448 306342 327500 306348
rect 327460 293282 327488 306342
rect 327644 302234 327672 310406
rect 327920 306474 327948 310420
rect 327908 306468 327960 306474
rect 327908 306410 327960 306416
rect 328104 306406 328132 310420
rect 328196 310406 328394 310434
rect 328196 306542 328224 310406
rect 328184 306536 328236 306542
rect 328184 306478 328236 306484
rect 328092 306400 328144 306406
rect 328092 306342 328144 306348
rect 328460 306400 328512 306406
rect 328460 306342 328512 306348
rect 328564 306354 328592 310420
rect 328762 310406 328960 310434
rect 327644 302206 327764 302234
rect 327736 296714 327764 302206
rect 327552 296686 327764 296714
rect 327552 294710 327580 296686
rect 327540 294704 327592 294710
rect 327540 294646 327592 294652
rect 327448 293276 327500 293282
rect 327448 293218 327500 293224
rect 327356 275324 327408 275330
rect 327356 275266 327408 275272
rect 327264 269884 327316 269890
rect 327264 269826 327316 269832
rect 328472 268462 328500 306342
rect 328564 306326 328868 306354
rect 328644 305380 328696 305386
rect 328644 305322 328696 305328
rect 328552 305244 328604 305250
rect 328552 305186 328604 305192
rect 328564 271182 328592 305186
rect 328656 274038 328684 305322
rect 328736 305312 328788 305318
rect 328736 305254 328788 305260
rect 328748 291854 328776 305254
rect 328840 294642 328868 306326
rect 328932 301578 328960 310406
rect 329024 305386 329052 310420
rect 329208 306406 329236 310420
rect 329196 306400 329248 306406
rect 329196 306342 329248 306348
rect 329012 305380 329064 305386
rect 329012 305322 329064 305328
rect 329392 305318 329420 310420
rect 329484 310406 329682 310434
rect 329380 305312 329432 305318
rect 329380 305254 329432 305260
rect 329484 305250 329512 310406
rect 329852 306474 329880 310420
rect 329944 310406 330142 310434
rect 329840 306468 329892 306474
rect 329840 306410 329892 306416
rect 329944 306354 329972 310406
rect 330312 306354 330340 310420
rect 329852 306326 329972 306354
rect 330036 306326 330340 306354
rect 329472 305244 329524 305250
rect 329472 305186 329524 305192
rect 328920 301572 328972 301578
rect 328920 301514 328972 301520
rect 328828 294636 328880 294642
rect 328828 294578 328880 294584
rect 328736 291848 328788 291854
rect 328736 291790 328788 291796
rect 328644 274032 328696 274038
rect 328644 273974 328696 273980
rect 328552 271176 328604 271182
rect 328552 271118 328604 271124
rect 328460 268456 328512 268462
rect 328460 268398 328512 268404
rect 327172 246492 327224 246498
rect 327172 246434 327224 246440
rect 329852 246430 329880 306326
rect 329932 305244 329984 305250
rect 329932 305186 329984 305192
rect 329944 247722 329972 305186
rect 330036 250510 330064 306326
rect 330208 305380 330260 305386
rect 330208 305322 330260 305328
rect 330116 305312 330168 305318
rect 330116 305254 330168 305260
rect 330128 254590 330156 305254
rect 330220 260166 330248 305322
rect 330496 302234 330524 310420
rect 330588 310406 330786 310434
rect 330588 305250 330616 310406
rect 330668 306468 330720 306474
rect 330668 306410 330720 306416
rect 330576 305244 330628 305250
rect 330576 305186 330628 305192
rect 330680 302234 330708 306410
rect 330956 305318 330984 310420
rect 331140 305386 331168 310420
rect 331220 306536 331272 306542
rect 331220 306478 331272 306484
rect 331128 305380 331180 305386
rect 331128 305322 331180 305328
rect 330944 305312 330996 305318
rect 330944 305254 330996 305260
rect 330312 302206 330524 302234
rect 330588 302206 330708 302234
rect 330312 261526 330340 302206
rect 330588 296714 330616 302206
rect 330404 296686 330616 296714
rect 330404 278050 330432 296686
rect 330392 278044 330444 278050
rect 330392 277986 330444 277992
rect 330300 261520 330352 261526
rect 330300 261462 330352 261468
rect 330208 260160 330260 260166
rect 330208 260102 330260 260108
rect 330116 254584 330168 254590
rect 330116 254526 330168 254532
rect 330024 250504 330076 250510
rect 330024 250446 330076 250452
rect 329932 247716 329984 247722
rect 329932 247658 329984 247664
rect 329840 246424 329892 246430
rect 329840 246366 329892 246372
rect 331232 246362 331260 306478
rect 331312 306332 331364 306338
rect 331312 306274 331364 306280
rect 331324 265742 331352 306274
rect 331416 305561 331444 310420
rect 331600 306354 331628 310420
rect 331784 306542 331812 310420
rect 331876 310406 332074 310434
rect 331772 306536 331824 306542
rect 331772 306478 331824 306484
rect 331508 306326 331628 306354
rect 331402 305552 331458 305561
rect 331402 305487 331458 305496
rect 331404 305380 331456 305386
rect 331404 305322 331456 305328
rect 331416 268394 331444 305322
rect 331508 269822 331536 306326
rect 331876 306252 331904 310406
rect 331956 306468 332008 306474
rect 331956 306410 332008 306416
rect 331600 306224 331904 306252
rect 331600 289202 331628 306224
rect 331678 305552 331734 305561
rect 331678 305487 331734 305496
rect 331692 290562 331720 305487
rect 331968 305318 331996 306410
rect 332244 305386 332272 310420
rect 332336 310406 332534 310434
rect 332336 306338 332364 310406
rect 332704 306474 332732 310420
rect 332692 306468 332744 306474
rect 332692 306410 332744 306416
rect 332888 306354 332916 310420
rect 332324 306332 332376 306338
rect 332324 306274 332376 306280
rect 332600 306332 332652 306338
rect 332600 306274 332652 306280
rect 332704 306326 332916 306354
rect 332980 310406 333178 310434
rect 332508 305584 332560 305590
rect 332508 305526 332560 305532
rect 332520 305454 332548 305526
rect 332508 305448 332560 305454
rect 332508 305390 332560 305396
rect 332232 305380 332284 305386
rect 332232 305322 332284 305328
rect 331956 305312 332008 305318
rect 331956 305254 332008 305260
rect 331680 290556 331732 290562
rect 331680 290498 331732 290504
rect 331588 289196 331640 289202
rect 331588 289138 331640 289144
rect 331496 269816 331548 269822
rect 331496 269758 331548 269764
rect 331404 268388 331456 268394
rect 331404 268330 331456 268336
rect 331312 265736 331364 265742
rect 331312 265678 331364 265684
rect 332612 251870 332640 306274
rect 332704 267034 332732 306326
rect 332876 305584 332928 305590
rect 332876 305526 332928 305532
rect 332784 305380 332836 305386
rect 332784 305322 332836 305328
rect 332796 272542 332824 305322
rect 332888 287706 332916 305526
rect 332980 297498 333008 310406
rect 333060 306468 333112 306474
rect 333060 306410 333112 306416
rect 333072 298790 333100 306410
rect 333348 305590 333376 310420
rect 333336 305584 333388 305590
rect 333336 305526 333388 305532
rect 333532 305386 333560 310420
rect 333624 310406 333822 310434
rect 333624 306338 333652 310406
rect 333992 306542 334020 310420
rect 334190 310406 334296 310434
rect 334268 307902 334296 310406
rect 334256 307896 334308 307902
rect 334256 307838 334308 307844
rect 333980 306536 334032 306542
rect 333980 306478 334032 306484
rect 333980 306400 334032 306406
rect 333980 306342 334032 306348
rect 333612 306332 333664 306338
rect 333612 306274 333664 306280
rect 333520 305380 333572 305386
rect 333520 305322 333572 305328
rect 333060 298784 333112 298790
rect 333060 298726 333112 298732
rect 332968 297492 333020 297498
rect 332968 297434 333020 297440
rect 332876 287700 332928 287706
rect 332876 287642 332928 287648
rect 333992 283626 334020 306342
rect 334072 306332 334124 306338
rect 334072 306274 334124 306280
rect 334084 289134 334112 306274
rect 334452 305674 334480 310420
rect 334636 307222 334664 310420
rect 334728 310406 334926 310434
rect 334624 307216 334676 307222
rect 334624 307158 334676 307164
rect 334532 306536 334584 306542
rect 334532 306478 334584 306484
rect 334176 305646 334480 305674
rect 334176 290494 334204 305646
rect 334256 305584 334308 305590
rect 334256 305526 334308 305532
rect 334268 297430 334296 305526
rect 334544 304298 334572 306478
rect 334728 306338 334756 310406
rect 334808 307896 334860 307902
rect 334808 307838 334860 307844
rect 334716 306332 334768 306338
rect 334716 306274 334768 306280
rect 334532 304292 334584 304298
rect 334532 304234 334584 304240
rect 334820 301510 334848 307838
rect 335096 306406 335124 310420
rect 335084 306400 335136 306406
rect 335084 306342 335136 306348
rect 335280 305590 335308 310420
rect 335372 310406 335570 310434
rect 335268 305584 335320 305590
rect 335268 305526 335320 305532
rect 334808 301504 334860 301510
rect 334808 301446 334860 301452
rect 334256 297424 334308 297430
rect 334256 297366 334308 297372
rect 334164 290488 334216 290494
rect 334164 290430 334216 290436
rect 334072 289128 334124 289134
rect 334072 289070 334124 289076
rect 333980 283620 334032 283626
rect 333980 283562 334032 283568
rect 332784 272536 332836 272542
rect 332784 272478 332836 272484
rect 332692 267028 332744 267034
rect 332692 266970 332744 266976
rect 332600 251864 332652 251870
rect 332600 251806 332652 251812
rect 335372 249082 335400 310406
rect 335740 306490 335768 310420
rect 335464 306462 335768 306490
rect 335464 253298 335492 306462
rect 335636 306400 335688 306406
rect 335636 306342 335688 306348
rect 335544 305584 335596 305590
rect 335544 305526 335596 305532
rect 335452 253292 335504 253298
rect 335452 253234 335504 253240
rect 335556 253230 335584 305526
rect 335648 253366 335676 306342
rect 335728 306332 335780 306338
rect 335728 306274 335780 306280
rect 335740 265674 335768 306274
rect 335924 296714 335952 310420
rect 336016 310406 336214 310434
rect 336016 306338 336044 310406
rect 336004 306332 336056 306338
rect 336004 306274 336056 306280
rect 336384 305590 336412 310420
rect 336568 306406 336596 310420
rect 336556 306400 336608 306406
rect 336556 306342 336608 306348
rect 336372 305584 336424 305590
rect 336372 305526 336424 305532
rect 335832 296686 335952 296714
rect 335832 286346 335860 296686
rect 335820 286340 335872 286346
rect 335820 286282 335872 286288
rect 336844 273970 336872 310420
rect 336924 306332 336976 306338
rect 336924 306274 336976 306280
rect 336936 300830 336964 306274
rect 336924 300824 336976 300830
rect 336924 300766 336976 300772
rect 336832 273964 336884 273970
rect 336832 273906 336884 273912
rect 335728 265668 335780 265674
rect 335728 265610 335780 265616
rect 335636 253360 335688 253366
rect 335636 253302 335688 253308
rect 335544 253224 335596 253230
rect 335544 253166 335596 253172
rect 335360 249076 335412 249082
rect 335360 249018 335412 249024
rect 331220 246356 331272 246362
rect 331220 246298 331272 246304
rect 306380 244870 306432 244876
rect 327078 244896 327134 244905
rect 327078 244831 327134 244840
rect 301042 244760 301098 244769
rect 337028 244730 337056 310420
rect 337120 310406 337318 310434
rect 337120 306338 337148 310406
rect 337488 308310 337516 310420
rect 337476 308304 337528 308310
rect 337476 308246 337528 308252
rect 337672 308174 337700 310420
rect 337948 308417 337976 310420
rect 337934 308408 337990 308417
rect 337934 308343 337990 308352
rect 337660 308168 337712 308174
rect 337660 308110 337712 308116
rect 337108 306332 337160 306338
rect 337108 306274 337160 306280
rect 338132 302734 338160 310420
rect 338212 306332 338264 306338
rect 338212 306274 338264 306280
rect 338120 302728 338172 302734
rect 338120 302670 338172 302676
rect 338224 300082 338252 306274
rect 338316 300762 338344 310420
rect 338592 309126 338620 310420
rect 338580 309120 338632 309126
rect 338580 309062 338632 309068
rect 338776 305454 338804 310420
rect 338960 306241 338988 310420
rect 339052 310406 339250 310434
rect 338946 306232 339002 306241
rect 338946 306167 339002 306176
rect 338764 305448 338816 305454
rect 338764 305390 338816 305396
rect 339052 302234 339080 310406
rect 339420 306338 339448 310420
rect 339696 306354 339724 310420
rect 339408 306332 339460 306338
rect 339408 306274 339460 306280
rect 339592 306332 339644 306338
rect 339696 306326 339816 306354
rect 339592 306274 339644 306280
rect 338408 302206 339080 302234
rect 338304 300756 338356 300762
rect 338304 300698 338356 300704
rect 338212 300076 338264 300082
rect 338212 300018 338264 300024
rect 338408 297838 338436 302206
rect 338396 297832 338448 297838
rect 338396 297774 338448 297780
rect 339604 247586 339632 306274
rect 339684 305584 339736 305590
rect 339684 305526 339736 305532
rect 339696 297702 339724 305526
rect 339684 297696 339736 297702
rect 339684 297638 339736 297644
rect 339592 247580 339644 247586
rect 339592 247522 339644 247528
rect 339788 244798 339816 306326
rect 339880 305318 339908 310420
rect 339868 305312 339920 305318
rect 339868 305254 339920 305260
rect 340064 303385 340092 310420
rect 340156 310406 340354 310434
rect 340156 305590 340184 310406
rect 340144 305584 340196 305590
rect 340144 305526 340196 305532
rect 340050 303376 340106 303385
rect 340050 303311 340106 303320
rect 340524 300014 340552 310420
rect 340708 306338 340736 310420
rect 340880 308440 340932 308446
rect 340880 308382 340932 308388
rect 340696 306332 340748 306338
rect 340696 306274 340748 306280
rect 340892 305522 340920 308382
rect 340984 306270 341012 310420
rect 341168 308394 341196 310420
rect 341352 308394 341380 310420
rect 341076 308366 341196 308394
rect 341260 308366 341380 308394
rect 341444 310406 341642 310434
rect 340972 306264 341024 306270
rect 340972 306206 341024 306212
rect 340880 305516 340932 305522
rect 340880 305458 340932 305464
rect 341076 303249 341104 308366
rect 341156 308304 341208 308310
rect 341156 308246 341208 308252
rect 341062 303240 341118 303249
rect 341062 303175 341118 303184
rect 340512 300008 340564 300014
rect 340512 299950 340564 299956
rect 341168 246294 341196 308246
rect 341260 303618 341288 308366
rect 341248 303612 341300 303618
rect 341248 303554 341300 303560
rect 341444 299946 341472 310406
rect 341812 308310 341840 310420
rect 341904 310406 342102 310434
rect 341904 308446 341932 310406
rect 342168 309120 342220 309126
rect 342168 309062 342220 309068
rect 341892 308440 341944 308446
rect 341892 308382 341944 308388
rect 341800 308304 341852 308310
rect 342180 308292 342208 309062
rect 342272 308394 342300 310420
rect 342470 310406 342668 310434
rect 342536 308440 342588 308446
rect 342272 308366 342484 308394
rect 342640 308428 342668 310406
rect 342732 308666 342760 310420
rect 342916 309126 342944 310420
rect 342904 309120 342956 309126
rect 342904 309062 342956 309068
rect 342732 308638 343036 308666
rect 342640 308400 342852 308428
rect 342536 308382 342588 308388
rect 342180 308264 342300 308292
rect 341800 308246 341852 308252
rect 342272 306202 342300 308264
rect 342352 308236 342404 308242
rect 342352 308178 342404 308184
rect 342260 306196 342312 306202
rect 342260 306138 342312 306144
rect 342364 303550 342392 308178
rect 342352 303544 342404 303550
rect 342352 303486 342404 303492
rect 342456 303113 342484 308366
rect 342442 303104 342498 303113
rect 342442 303039 342498 303048
rect 342548 302802 342576 308382
rect 342628 308304 342680 308310
rect 342628 308246 342680 308252
rect 342536 302796 342588 302802
rect 342536 302738 342588 302744
rect 341432 299940 341484 299946
rect 341432 299882 341484 299888
rect 341156 246288 341208 246294
rect 341156 246230 341208 246236
rect 342640 244866 342668 308246
rect 342824 302870 342852 308400
rect 342812 302864 342864 302870
rect 342812 302806 342864 302812
rect 343008 296714 343036 308638
rect 343100 308242 343128 310420
rect 343192 310406 343390 310434
rect 343192 308446 343220 310406
rect 343180 308440 343232 308446
rect 343180 308382 343232 308388
rect 343560 308310 343588 310420
rect 343744 309346 343772 310420
rect 343652 309318 343772 309346
rect 343836 310406 344034 310434
rect 343652 308446 343680 309318
rect 343836 308802 343864 310406
rect 343744 308774 343864 308802
rect 343640 308440 343692 308446
rect 343640 308382 343692 308388
rect 343548 308304 343600 308310
rect 343548 308246 343600 308252
rect 343088 308236 343140 308242
rect 343088 308178 343140 308184
rect 343640 307284 343692 307290
rect 343640 307226 343692 307232
rect 343652 305454 343680 307226
rect 343640 305448 343692 305454
rect 343640 305390 343692 305396
rect 343744 303482 343772 308774
rect 344204 308666 344232 310420
rect 343836 308638 344232 308666
rect 344296 310406 344494 310434
rect 343732 303476 343784 303482
rect 343732 303418 343784 303424
rect 343836 297770 343864 308638
rect 343916 308440 343968 308446
rect 344296 308394 344324 310406
rect 343916 308382 343968 308388
rect 343824 297764 343876 297770
rect 343824 297706 343876 297712
rect 342732 296686 343036 296714
rect 342732 247042 342760 296686
rect 342720 247036 342772 247042
rect 342720 246978 342772 246984
rect 342628 244860 342680 244866
rect 342628 244802 342680 244808
rect 339776 244792 339828 244798
rect 339776 244734 339828 244740
rect 301042 244695 301098 244704
rect 337016 244724 337068 244730
rect 337016 244666 337068 244672
rect 300768 243772 300820 243778
rect 300768 243714 300820 243720
rect 343928 243710 343956 308382
rect 344020 308366 344324 308394
rect 344020 252074 344048 308366
rect 344664 307290 344692 310420
rect 344652 307284 344704 307290
rect 344652 307226 344704 307232
rect 344848 303414 344876 310420
rect 345032 310406 345138 310434
rect 344836 303408 344888 303414
rect 344836 303350 344888 303356
rect 345032 300694 345060 310406
rect 345204 308440 345256 308446
rect 345204 308382 345256 308388
rect 345112 308372 345164 308378
rect 345112 308314 345164 308320
rect 345124 303278 345152 308314
rect 345112 303272 345164 303278
rect 345112 303214 345164 303220
rect 345020 300688 345072 300694
rect 345020 300630 345072 300636
rect 344008 252068 344060 252074
rect 344008 252010 344060 252016
rect 345216 248334 345244 308382
rect 345308 308310 345336 310420
rect 345492 308394 345520 310420
rect 345400 308366 345520 308394
rect 345584 310406 345782 310434
rect 345584 308378 345612 310406
rect 345952 308446 345980 310420
rect 345940 308440 345992 308446
rect 345940 308382 345992 308388
rect 345572 308372 345624 308378
rect 345296 308304 345348 308310
rect 345296 308246 345348 308252
rect 345296 308168 345348 308174
rect 345296 308110 345348 308116
rect 345308 300490 345336 308110
rect 345296 300484 345348 300490
rect 345296 300426 345348 300432
rect 345204 248328 345256 248334
rect 345204 248270 345256 248276
rect 343916 243704 343968 243710
rect 343916 243646 343968 243652
rect 345400 243642 345428 308366
rect 345572 308314 345624 308320
rect 345480 308304 345532 308310
rect 345480 308246 345532 308252
rect 345492 246974 345520 308246
rect 346136 308174 346164 310420
rect 346124 308168 346176 308174
rect 346124 308110 346176 308116
rect 346412 303210 346440 310420
rect 346610 310406 346808 310434
rect 346584 308440 346636 308446
rect 346584 308382 346636 308388
rect 346400 303204 346452 303210
rect 346400 303146 346452 303152
rect 346596 300626 346624 308382
rect 346676 308372 346728 308378
rect 346676 308314 346728 308320
rect 346584 300620 346636 300626
rect 346584 300562 346636 300568
rect 346688 248198 346716 308314
rect 346676 248192 346728 248198
rect 346676 248134 346728 248140
rect 346780 247654 346808 310406
rect 346872 308446 346900 310420
rect 347056 308689 347084 310420
rect 347042 308680 347098 308689
rect 347042 308615 347098 308624
rect 346860 308440 346912 308446
rect 346860 308382 346912 308388
rect 347240 308378 347268 310420
rect 347332 310406 347530 310434
rect 347228 308372 347280 308378
rect 347228 308314 347280 308320
rect 347332 300422 347360 310406
rect 347700 308582 347728 310420
rect 347898 310406 348004 310434
rect 347688 308576 347740 308582
rect 347688 308518 347740 308524
rect 347320 300416 347372 300422
rect 347320 300358 347372 300364
rect 347976 248402 348004 310406
rect 348160 308922 348188 310420
rect 348344 308961 348372 310420
rect 348330 308952 348386 308961
rect 348148 308916 348200 308922
rect 348330 308887 348386 308896
rect 348148 308858 348200 308864
rect 348528 296714 348556 310420
rect 348804 308718 348832 310420
rect 348792 308712 348844 308718
rect 348792 308654 348844 308660
rect 348988 308514 349016 310420
rect 348976 308508 349028 308514
rect 348976 308450 349028 308456
rect 348252 296686 348556 296714
rect 347964 248396 348016 248402
rect 347964 248338 348016 248344
rect 348252 248130 348280 296686
rect 348240 248124 348292 248130
rect 348240 248066 348292 248072
rect 346768 247648 346820 247654
rect 346768 247590 346820 247596
rect 345480 246968 345532 246974
rect 345480 246910 345532 246916
rect 349264 246702 349292 310420
rect 349448 308650 349476 310420
rect 349632 308825 349660 310420
rect 349724 310406 349922 310434
rect 349618 308816 349674 308825
rect 349618 308751 349674 308760
rect 349436 308644 349488 308650
rect 349436 308586 349488 308592
rect 349344 308440 349396 308446
rect 349344 308382 349396 308388
rect 349356 300218 349384 308382
rect 349344 300212 349396 300218
rect 349344 300154 349396 300160
rect 349724 296714 349752 310406
rect 350092 308446 350120 310420
rect 350080 308440 350132 308446
rect 350080 308382 350132 308388
rect 350276 308242 350304 310420
rect 350552 308258 350580 310420
rect 350736 308632 350764 310420
rect 350920 308990 350948 310420
rect 350908 308984 350960 308990
rect 350908 308926 350960 308932
rect 350736 308604 351132 308632
rect 350264 308236 350316 308242
rect 350552 308230 350948 308258
rect 350264 308178 350316 308184
rect 350816 308168 350868 308174
rect 350816 308110 350868 308116
rect 350632 308100 350684 308106
rect 350632 308042 350684 308048
rect 350644 306134 350672 308042
rect 350724 306604 350776 306610
rect 350724 306546 350776 306552
rect 350632 306128 350684 306134
rect 350632 306070 350684 306076
rect 349448 296686 349752 296714
rect 349448 246838 349476 296686
rect 350736 248266 350764 306546
rect 350828 267170 350856 308110
rect 350816 267164 350868 267170
rect 350816 267106 350868 267112
rect 350724 248260 350776 248266
rect 350724 248202 350776 248208
rect 349436 246832 349488 246838
rect 349436 246774 349488 246780
rect 350920 246770 350948 308230
rect 351104 300354 351132 308604
rect 351092 300348 351144 300354
rect 351092 300290 351144 300296
rect 351196 296714 351224 310420
rect 351380 308106 351408 310420
rect 351472 310406 351670 310434
rect 351472 308174 351500 310406
rect 351460 308168 351512 308174
rect 351460 308110 351512 308116
rect 351368 308100 351420 308106
rect 351368 308042 351420 308048
rect 351840 306610 351868 310420
rect 352024 308854 352052 310420
rect 352012 308848 352064 308854
rect 352012 308790 352064 308796
rect 352300 308553 352328 310420
rect 352286 308544 352342 308553
rect 352286 308479 352342 308488
rect 352484 308446 352512 310420
rect 352472 308440 352524 308446
rect 352472 308382 352524 308388
rect 351828 306604 351880 306610
rect 351828 306546 351880 306552
rect 352668 300665 352696 310420
rect 352944 309058 352972 310420
rect 352932 309052 352984 309058
rect 352932 308994 352984 309000
rect 353128 308514 353156 310420
rect 353404 310406 353602 310434
rect 353116 308508 353168 308514
rect 353116 308450 353168 308456
rect 353404 306105 353432 310406
rect 353390 306096 353446 306105
rect 353390 306031 353446 306040
rect 353680 305726 353708 310490
rect 353772 308582 353800 310420
rect 354048 308786 354076 310420
rect 354036 308780 354088 308786
rect 354036 308722 354088 308728
rect 353760 308576 353812 308582
rect 353760 308518 353812 308524
rect 354232 305998 354260 310420
rect 354416 308718 354444 310420
rect 354404 308712 354456 308718
rect 354404 308654 354456 308660
rect 354692 308378 354720 310420
rect 354876 308530 354904 310420
rect 355060 308990 355088 310420
rect 355152 310406 355350 310434
rect 355048 308984 355100 308990
rect 355048 308926 355100 308932
rect 354784 308502 354904 308530
rect 354680 308372 354732 308378
rect 354680 308314 354732 308320
rect 354784 308258 354812 308502
rect 354864 308372 354916 308378
rect 354864 308314 354916 308320
rect 354692 308230 354812 308258
rect 354220 305992 354272 305998
rect 354220 305934 354272 305940
rect 354692 305930 354720 308230
rect 354772 308168 354824 308174
rect 354772 308110 354824 308116
rect 354680 305924 354732 305930
rect 354680 305866 354732 305872
rect 354784 305862 354812 308110
rect 354876 306066 354904 308314
rect 354864 306060 354916 306066
rect 354864 306002 354916 306008
rect 354772 305856 354824 305862
rect 354772 305798 354824 305804
rect 353668 305720 353720 305726
rect 353668 305662 353720 305668
rect 355152 303346 355180 310406
rect 355520 308174 355548 310420
rect 355704 308786 355732 310420
rect 355796 310406 355994 310434
rect 355692 308780 355744 308786
rect 355692 308722 355744 308728
rect 355508 308168 355560 308174
rect 355508 308110 355560 308116
rect 355140 303340 355192 303346
rect 355140 303282 355192 303288
rect 352654 300656 352710 300665
rect 352654 300591 352710 300600
rect 355796 300393 355824 310406
rect 356244 308644 356296 308650
rect 356244 308586 356296 308592
rect 356152 308372 356204 308378
rect 356152 308314 356204 308320
rect 356060 308304 356112 308310
rect 356060 308246 356112 308252
rect 355782 300384 355838 300393
rect 355782 300319 355838 300328
rect 351012 296686 351224 296714
rect 351012 246906 351040 296686
rect 351000 246900 351052 246906
rect 351000 246842 351052 246848
rect 350908 246764 350960 246770
rect 350908 246706 350960 246712
rect 349252 246696 349304 246702
rect 349252 246638 349304 246644
rect 345388 243636 345440 243642
rect 345388 243578 345440 243584
rect 356072 243574 356100 308246
rect 356164 305794 356192 308314
rect 356152 305788 356204 305794
rect 356152 305730 356204 305736
rect 356256 248334 356284 308586
rect 356348 250782 356376 310542
rect 356440 308650 356468 310420
rect 356428 308644 356480 308650
rect 356428 308586 356480 308592
rect 356624 308394 356652 310420
rect 356440 308366 356652 308394
rect 356808 308378 356836 310420
rect 356900 310406 357098 310434
rect 356796 308372 356848 308378
rect 356440 300529 356468 308366
rect 356796 308314 356848 308320
rect 356426 300520 356482 300529
rect 356426 300455 356482 300464
rect 356900 296714 356928 310406
rect 357268 308310 357296 310420
rect 357256 308304 357308 308310
rect 357256 308246 357308 308252
rect 357452 305658 357480 310420
rect 357728 308394 357756 310420
rect 357532 308372 357584 308378
rect 357728 308366 357848 308394
rect 357532 308314 357584 308320
rect 357440 305652 357492 305658
rect 357440 305594 357492 305600
rect 357544 303142 357572 308314
rect 357716 308304 357768 308310
rect 357716 308246 357768 308252
rect 357624 308236 357676 308242
rect 357624 308178 357676 308184
rect 357532 303136 357584 303142
rect 357532 303078 357584 303084
rect 357636 300558 357664 308178
rect 357624 300552 357676 300558
rect 357624 300494 357676 300500
rect 356532 296686 356928 296714
rect 356336 250776 356388 250782
rect 356336 250718 356388 250724
rect 356244 248328 356296 248334
rect 356244 248270 356296 248276
rect 356532 244866 356560 296686
rect 357728 248130 357756 308246
rect 357820 248198 357848 308366
rect 357912 300286 357940 310420
rect 358096 308378 358124 310420
rect 358188 310406 358386 310434
rect 358084 308372 358136 308378
rect 358084 308314 358136 308320
rect 358188 308310 358216 310406
rect 358176 308304 358228 308310
rect 358176 308246 358228 308252
rect 358556 308242 358584 310420
rect 358832 308394 358860 310420
rect 359016 308650 359044 310420
rect 359004 308644 359056 308650
rect 359004 308586 359056 308592
rect 359200 308394 359228 310420
rect 359280 308644 359332 308650
rect 359280 308586 359332 308592
rect 358832 308366 358952 308394
rect 358544 308236 358596 308242
rect 358544 308178 358596 308184
rect 358820 308168 358872 308174
rect 358820 308110 358872 308116
rect 358832 303006 358860 308110
rect 358924 303074 358952 308366
rect 359016 308366 359228 308394
rect 358912 303068 358964 303074
rect 358912 303010 358964 303016
rect 358820 303000 358872 303006
rect 358820 302942 358872 302948
rect 357900 300280 357952 300286
rect 357900 300222 357952 300228
rect 359016 297634 359044 308366
rect 359188 308304 359240 308310
rect 359188 308246 359240 308252
rect 359096 308236 359148 308242
rect 359096 308178 359148 308184
rect 359108 302938 359136 308178
rect 359096 302932 359148 302938
rect 359096 302874 359148 302880
rect 359200 300257 359228 308246
rect 359292 308106 359320 308586
rect 359476 308174 359504 310420
rect 359464 308168 359516 308174
rect 359464 308110 359516 308116
rect 359280 308100 359332 308106
rect 359280 308042 359332 308048
rect 359660 307986 359688 310420
rect 359844 308310 359872 310420
rect 359936 310406 360134 310434
rect 359832 308304 359884 308310
rect 359832 308246 359884 308252
rect 359936 308242 359964 310406
rect 360304 308802 360332 310420
rect 360120 308774 360332 308802
rect 360120 308394 360148 308774
rect 360120 308366 360332 308394
rect 360200 308304 360252 308310
rect 360200 308246 360252 308252
rect 359924 308236 359976 308242
rect 359924 308178 359976 308184
rect 359292 307958 359688 307986
rect 359186 300248 359242 300257
rect 359186 300183 359242 300192
rect 359004 297628 359056 297634
rect 359004 297570 359056 297576
rect 359292 248266 359320 307958
rect 359372 307896 359424 307902
rect 359372 307838 359424 307844
rect 359384 250782 359412 307838
rect 360212 300150 360240 308246
rect 360200 300144 360252 300150
rect 360200 300086 360252 300092
rect 359372 250776 359424 250782
rect 359372 250718 359424 250724
rect 360304 248402 360332 308366
rect 360488 308310 360516 310420
rect 360580 310406 360778 310434
rect 360476 308304 360528 308310
rect 360476 308246 360528 308252
rect 360580 308122 360608 310406
rect 360396 308094 360608 308122
rect 360396 263090 360424 308094
rect 360948 296714 360976 310420
rect 361132 309806 361160 443006
rect 362236 325650 362264 446354
rect 363604 446344 363656 446350
rect 363604 446286 363656 446292
rect 362316 446276 362368 446282
rect 362316 446218 362368 446224
rect 362328 439550 362356 446218
rect 362316 439544 362368 439550
rect 362316 439486 362368 439492
rect 362224 325644 362276 325650
rect 362224 325586 362276 325592
rect 361120 309800 361172 309806
rect 361120 309742 361172 309748
rect 360488 296686 360976 296714
rect 360384 263084 360436 263090
rect 360384 263026 360436 263032
rect 360292 248396 360344 248402
rect 360292 248338 360344 248344
rect 359280 248260 359332 248266
rect 359280 248202 359332 248208
rect 357808 248192 357860 248198
rect 357808 248134 357860 248140
rect 357716 248124 357768 248130
rect 357716 248066 357768 248072
rect 356520 244860 356572 244866
rect 356520 244802 356572 244808
rect 360488 244798 360516 296686
rect 363616 258738 363644 446286
rect 364996 260234 365024 446422
rect 373264 446208 373316 446214
rect 373264 446150 373316 446156
rect 369124 443692 369176 443698
rect 369124 443634 369176 443640
rect 367744 443624 367796 443630
rect 367744 443566 367796 443572
rect 367756 273222 367784 443566
rect 369136 379506 369164 443634
rect 369124 379500 369176 379506
rect 369124 379442 369176 379448
rect 367744 273216 367796 273222
rect 367744 273158 367796 273164
rect 364984 260228 365036 260234
rect 364984 260170 365036 260176
rect 363604 258732 363656 258738
rect 363604 258674 363656 258680
rect 373276 257378 373304 446150
rect 458824 445868 458876 445874
rect 458824 445810 458876 445816
rect 446404 443216 446456 443222
rect 446404 443158 446456 443164
rect 438032 308780 438084 308786
rect 438032 308722 438084 308728
rect 436836 308712 436888 308718
rect 436836 308654 436888 308660
rect 436744 264444 436796 264450
rect 436744 264386 436796 264392
rect 373264 257372 373316 257378
rect 373264 257314 373316 257320
rect 360476 244792 360528 244798
rect 360476 244734 360528 244740
rect 356060 243568 356112 243574
rect 356060 243510 356112 243516
rect 348238 159896 348294 159905
rect 348238 159831 348294 159840
rect 350998 159896 351054 159905
rect 350998 159831 351054 159840
rect 356058 159896 356114 159905
rect 356058 159831 356114 159840
rect 358450 159896 358506 159905
rect 358450 159831 358506 159840
rect 360934 159896 360990 159905
rect 360934 159831 360990 159840
rect 368294 159896 368350 159905
rect 368294 159831 368350 159840
rect 299480 159656 299532 159662
rect 299480 159598 299532 159604
rect 299388 159112 299440 159118
rect 299388 159054 299440 159060
rect 299308 158902 299428 158930
rect 299204 158296 299256 158302
rect 299204 158238 299256 158244
rect 299400 158234 299428 158902
rect 299388 158228 299440 158234
rect 299388 158170 299440 158176
rect 299400 157622 299428 158170
rect 299388 157616 299440 157622
rect 299388 157558 299440 157564
rect 299388 155372 299440 155378
rect 299388 155314 299440 155320
rect 299400 154970 299428 155314
rect 299388 154964 299440 154970
rect 299388 154906 299440 154912
rect 299112 152516 299164 152522
rect 299112 152458 299164 152464
rect 299020 8968 299072 8974
rect 299020 8910 299072 8916
rect 298100 7608 298152 7614
rect 298100 7550 298152 7556
rect 295524 6792 295576 6798
rect 295524 6734 295576 6740
rect 297272 4888 297324 4894
rect 297272 4830 297324 4836
rect 295432 4004 295484 4010
rect 295432 3946 295484 3952
rect 295248 3936 295300 3942
rect 295248 3878 295300 3884
rect 295156 3800 295208 3806
rect 295156 3742 295208 3748
rect 295064 3528 295116 3534
rect 295064 3470 295116 3476
rect 296076 3188 296128 3194
rect 296076 3130 296128 3136
rect 296088 480 296116 3130
rect 297284 480 297312 4830
rect 298468 4820 298520 4826
rect 298468 4762 298520 4768
rect 298480 480 298508 4762
rect 299492 3482 299520 159598
rect 309140 159588 309192 159594
rect 309140 159530 309192 159536
rect 302240 156528 302292 156534
rect 302240 156470 302292 156476
rect 300858 152416 300914 152425
rect 300858 152351 300914 152360
rect 299572 151224 299624 151230
rect 299572 151166 299624 151172
rect 299584 4214 299612 151166
rect 300872 16574 300900 152351
rect 302252 16574 302280 156470
rect 306380 155168 306432 155174
rect 306380 155110 306432 155116
rect 303620 149864 303672 149870
rect 303620 149806 303672 149812
rect 303632 16574 303660 149806
rect 305000 141500 305052 141506
rect 305000 141442 305052 141448
rect 305012 16574 305040 141442
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299572 4208 299624 4214
rect 299572 4150 299624 4156
rect 300768 4208 300820 4214
rect 300768 4150 300820 4156
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 4150
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 155110
rect 309152 16574 309180 159530
rect 327172 159520 327224 159526
rect 327172 159462 327224 159468
rect 316038 158672 316094 158681
rect 316038 158607 316094 158616
rect 317050 158672 317106 158681
rect 317050 158607 317106 158616
rect 319442 158672 319498 158681
rect 319442 158607 319498 158616
rect 320546 158672 320602 158681
rect 320546 158607 320602 158616
rect 321650 158672 321706 158681
rect 321650 158607 321706 158616
rect 323122 158672 323178 158681
rect 323122 158607 323178 158616
rect 316052 156874 316080 158607
rect 316040 156868 316092 156874
rect 316040 156810 316092 156816
rect 317064 156738 317092 158607
rect 319456 158098 319484 158607
rect 319444 158092 319496 158098
rect 319444 158034 319496 158040
rect 320560 157962 320588 158607
rect 320548 157956 320600 157962
rect 320548 157898 320600 157904
rect 321664 157894 321692 158607
rect 321652 157888 321704 157894
rect 321652 157830 321704 157836
rect 323136 156806 323164 158607
rect 324226 157856 324282 157865
rect 324226 157791 324282 157800
rect 323124 156800 323176 156806
rect 323124 156742 323176 156748
rect 317052 156732 317104 156738
rect 317052 156674 317104 156680
rect 313280 156596 313332 156602
rect 313280 156538 313332 156544
rect 310520 147008 310572 147014
rect 310520 146950 310572 146956
rect 310532 16574 310560 146950
rect 313292 16574 313320 156538
rect 324240 155446 324268 157791
rect 324870 157448 324926 157457
rect 324870 157383 324926 157392
rect 324228 155440 324280 155446
rect 324228 155382 324280 155388
rect 320180 155304 320232 155310
rect 320180 155246 320232 155252
rect 316040 153876 316092 153882
rect 316040 153818 316092 153824
rect 314660 145716 314712 145722
rect 314660 145658 314712 145664
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 313292 16546 313872 16574
rect 307944 13116 307996 13122
rect 307944 13058 307996 13064
rect 307956 480 307984 13058
rect 309048 6860 309100 6866
rect 309048 6802 309100 6808
rect 309060 480 309088 6802
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 312176 14476 312228 14482
rect 312176 14418 312228 14424
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 14418
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 145658
rect 316052 3398 316080 153818
rect 317420 144288 317472 144294
rect 317420 144230 317472 144236
rect 317432 16574 317460 144230
rect 318800 134564 318852 134570
rect 318800 134506 318852 134512
rect 318812 16574 318840 134506
rect 320192 16574 320220 155246
rect 324884 154222 324912 157383
rect 324872 154216 324924 154222
rect 324872 154158 324924 154164
rect 324320 152652 324372 152658
rect 324320 152594 324372 152600
rect 321560 142928 321612 142934
rect 321560 142870 321612 142876
rect 321572 16574 321600 142870
rect 322940 131776 322992 131782
rect 322940 131718 322992 131724
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316224 11756 316276 11762
rect 316224 11698 316276 11704
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 11698
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 131718
rect 324332 3210 324360 152594
rect 324412 151156 324464 151162
rect 324412 151098 324464 151104
rect 324424 3398 324452 151098
rect 325700 130416 325752 130422
rect 325700 130358 325752 130364
rect 325712 16574 325740 130358
rect 327184 16574 327212 159462
rect 338764 159452 338816 159458
rect 338764 159394 338816 159400
rect 338396 158704 338448 158710
rect 327538 158672 327594 158681
rect 327538 158607 327594 158616
rect 328274 158672 328330 158681
rect 328274 158607 328330 158616
rect 329930 158672 329986 158681
rect 329930 158607 329986 158616
rect 330298 158672 330354 158681
rect 330298 158607 330354 158616
rect 331218 158672 331274 158681
rect 331218 158607 331220 158616
rect 327552 158370 327580 158607
rect 328288 158506 328316 158607
rect 328276 158500 328328 158506
rect 328276 158442 328328 158448
rect 327540 158364 327592 158370
rect 327540 158306 327592 158312
rect 329944 158234 329972 158607
rect 329932 158228 329984 158234
rect 329932 158170 329984 158176
rect 329748 157480 329800 157486
rect 329748 157422 329800 157428
rect 327264 157412 327316 157418
rect 327264 157354 327316 157360
rect 327276 155378 327304 157354
rect 327264 155372 327316 155378
rect 327264 155314 327316 155320
rect 329760 154154 329788 157422
rect 330312 157078 330340 158607
rect 331272 158607 331274 158616
rect 332322 158672 332378 158681
rect 332322 158607 332378 158616
rect 333610 158672 333666 158681
rect 333610 158607 333666 158616
rect 334530 158672 334586 158681
rect 334530 158607 334586 158616
rect 335818 158672 335874 158681
rect 335818 158607 335874 158616
rect 336002 158672 336058 158681
rect 336002 158607 336058 158616
rect 336922 158672 336978 158681
rect 336922 158607 336978 158616
rect 338394 158672 338396 158681
rect 338448 158672 338450 158681
rect 338394 158607 338450 158616
rect 331220 158578 331272 158584
rect 332336 158302 332364 158607
rect 332324 158296 332376 158302
rect 332324 158238 332376 158244
rect 333624 158030 333652 158607
rect 333612 158024 333664 158030
rect 333612 157966 333664 157972
rect 331312 157548 331364 157554
rect 331312 157490 331364 157496
rect 330300 157072 330352 157078
rect 330300 157014 330352 157020
rect 331220 156664 331272 156670
rect 331220 156606 331272 156612
rect 329748 154148 329800 154154
rect 329748 154090 329800 154096
rect 328460 146940 328512 146946
rect 328460 146882 328512 146888
rect 328472 16574 328500 146882
rect 325712 16546 326384 16574
rect 327184 16546 328040 16574
rect 328472 16546 328776 16574
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330392 15904 330444 15910
rect 330392 15846 330444 15852
rect 330404 480 330432 15846
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 156606
rect 331324 154086 331352 157490
rect 334544 156942 334572 158607
rect 335832 157214 335860 158607
rect 336016 158166 336044 158607
rect 336004 158160 336056 158166
rect 336004 158102 336056 158108
rect 335820 157208 335872 157214
rect 335820 157150 335872 157156
rect 336936 157010 336964 158607
rect 338118 158264 338174 158273
rect 338118 158199 338174 158208
rect 336924 157004 336976 157010
rect 336924 156946 336976 156952
rect 334532 156936 334584 156942
rect 334532 156878 334584 156884
rect 338132 156398 338160 158199
rect 338120 156392 338172 156398
rect 338120 156334 338172 156340
rect 338120 155236 338172 155242
rect 338120 155178 338172 155184
rect 331312 154080 331364 154086
rect 331312 154022 331364 154028
rect 332600 148436 332652 148442
rect 332600 148378 332652 148384
rect 332612 3210 332640 148378
rect 335360 141432 335412 141438
rect 335360 141374 335412 141380
rect 332692 129056 332744 129062
rect 332692 128998 332744 129004
rect 332704 3398 332732 128998
rect 335372 16574 335400 141374
rect 336740 127628 336792 127634
rect 336740 127570 336792 127576
rect 336752 16574 336780 127570
rect 338132 16574 338160 155178
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 335084 4140 335136 4146
rect 335084 4082 335136 4088
rect 332692 3392 332744 3398
rect 332692 3334 332744 3340
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 332612 3182 332732 3210
rect 332704 480 332732 3182
rect 333900 480 333928 3334
rect 335096 480 335124 4082
rect 336292 480 336320 16546
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 338776 4146 338804 159394
rect 348252 159390 348280 159831
rect 348240 159384 348292 159390
rect 348240 159326 348292 159332
rect 351012 159322 351040 159831
rect 353574 159624 353630 159633
rect 353574 159559 353630 159568
rect 351000 159316 351052 159322
rect 351000 159258 351052 159264
rect 353588 159186 353616 159559
rect 356072 159254 356100 159831
rect 356060 159248 356112 159254
rect 356060 159190 356112 159196
rect 353576 159180 353628 159186
rect 353576 159122 353628 159128
rect 358464 158982 358492 159831
rect 358452 158976 358504 158982
rect 358452 158918 358504 158924
rect 360948 158914 360976 159831
rect 365902 159624 365958 159633
rect 365902 159559 365958 159568
rect 365916 159050 365944 159559
rect 368308 159118 368336 159831
rect 373998 159352 374054 159361
rect 373998 159287 374054 159296
rect 368296 159112 368348 159118
rect 368296 159054 368348 159060
rect 365904 159044 365956 159050
rect 365904 158986 365956 158992
rect 360936 158908 360988 158914
rect 360936 158850 360988 158856
rect 363420 158840 363472 158846
rect 363420 158782 363472 158788
rect 363432 158681 363460 158782
rect 370964 158772 371016 158778
rect 370964 158714 371016 158720
rect 370976 158681 371004 158714
rect 373448 158704 373500 158710
rect 339314 158672 339370 158681
rect 339314 158607 339370 158616
rect 340970 158672 341026 158681
rect 340970 158607 341026 158616
rect 343546 158672 343602 158681
rect 343546 158607 343602 158616
rect 347594 158672 347650 158681
rect 347594 158607 347650 158616
rect 354402 158672 354458 158681
rect 354402 158607 354458 158616
rect 355230 158672 355286 158681
rect 355230 158607 355286 158616
rect 356978 158672 357034 158681
rect 356978 158607 357034 158616
rect 363418 158672 363474 158681
rect 363418 158607 363474 158616
rect 370962 158672 371018 158681
rect 370962 158607 371018 158616
rect 373446 158672 373448 158681
rect 373500 158672 373502 158681
rect 373446 158607 373502 158616
rect 339328 157146 339356 158607
rect 340984 158574 341012 158607
rect 340972 158568 341024 158574
rect 340972 158510 341024 158516
rect 343560 158438 343588 158607
rect 343548 158432 343600 158438
rect 343548 158374 343600 158380
rect 343914 158264 343970 158273
rect 343914 158199 343970 158208
rect 341154 157992 341210 158001
rect 341154 157927 341210 157936
rect 339590 157856 339646 157865
rect 339590 157791 339646 157800
rect 339316 157140 339368 157146
rect 339316 157082 339368 157088
rect 339604 155582 339632 157791
rect 341168 155786 341196 157927
rect 342350 157856 342406 157865
rect 342350 157791 342406 157800
rect 341156 155780 341208 155786
rect 341156 155722 341208 155728
rect 342364 155650 342392 157791
rect 342352 155644 342404 155650
rect 342352 155586 342404 155592
rect 339592 155576 339644 155582
rect 339592 155518 339644 155524
rect 343928 155514 343956 158199
rect 345110 157992 345166 158001
rect 345110 157927 345166 157936
rect 346398 157992 346454 158001
rect 346398 157927 346454 157936
rect 345124 155922 345152 157927
rect 345754 157448 345810 157457
rect 345754 157383 345810 157392
rect 345112 155916 345164 155922
rect 345112 155858 345164 155864
rect 343916 155508 343968 155514
rect 343916 155450 343968 155456
rect 345768 154426 345796 157383
rect 346412 155854 346440 157927
rect 347608 157350 347636 158607
rect 348698 158264 348754 158273
rect 348698 158199 348754 158208
rect 353298 158264 353354 158273
rect 353298 158199 353354 158208
rect 347596 157344 347648 157350
rect 347596 157286 347648 157292
rect 346400 155848 346452 155854
rect 346400 155790 346452 155796
rect 348712 155718 348740 158199
rect 349802 157448 349858 157457
rect 349802 157383 349858 157392
rect 351090 157448 351146 157457
rect 351090 157383 351146 157392
rect 352194 157448 352250 157457
rect 352194 157383 352250 157392
rect 348700 155712 348752 155718
rect 348700 155654 348752 155660
rect 345756 154420 345808 154426
rect 345756 154362 345808 154368
rect 349816 154290 349844 157383
rect 351104 154562 351132 157383
rect 351092 154556 351144 154562
rect 351092 154498 351144 154504
rect 352208 154358 352236 157383
rect 353312 154494 353340 158199
rect 354416 157554 354444 158607
rect 354404 157548 354456 157554
rect 354404 157490 354456 157496
rect 355244 157418 355272 158607
rect 356992 157486 357020 158607
rect 356980 157480 357032 157486
rect 356980 157422 357032 157428
rect 355232 157412 355284 157418
rect 355232 157354 355284 157360
rect 353300 154488 353352 154494
rect 353300 154430 353352 154436
rect 352196 154352 352248 154358
rect 352196 154294 352248 154300
rect 349804 154284 349856 154290
rect 349804 154226 349856 154232
rect 349160 152584 349212 152590
rect 349160 152526 349212 152532
rect 340880 151088 340932 151094
rect 340880 151030 340932 151036
rect 339500 140072 339552 140078
rect 339500 140014 339552 140020
rect 338764 4140 338816 4146
rect 338764 4082 338816 4088
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 140014
rect 340892 3398 340920 151030
rect 345020 149796 345072 149802
rect 345020 149738 345072 149744
rect 342260 145648 342312 145654
rect 342260 145590 342312 145596
rect 340972 126268 341024 126274
rect 340972 126210 341024 126216
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 340984 480 341012 126210
rect 342272 16574 342300 145590
rect 343640 17264 343692 17270
rect 343640 17206 343692 17212
rect 343652 16574 343680 17206
rect 345032 16574 345060 149738
rect 346400 138712 346452 138718
rect 346400 138654 346452 138660
rect 346412 16574 346440 138654
rect 347780 29640 347832 29646
rect 347780 29582 347832 29588
rect 347792 16574 347820 29582
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3210 349200 152526
rect 357440 149728 357492 149734
rect 357440 149670 357492 149676
rect 351920 148368 351972 148374
rect 351920 148310 351972 148316
rect 350540 145580 350592 145586
rect 350540 145522 350592 145528
rect 349252 137284 349304 137290
rect 349252 137226 349304 137232
rect 349264 3398 349292 137226
rect 350552 16574 350580 145522
rect 351932 16574 351960 148310
rect 353300 144220 353352 144226
rect 353300 144162 353352 144168
rect 353312 16574 353340 144162
rect 354680 124908 354732 124914
rect 354680 124850 354732 124856
rect 354692 16574 354720 124850
rect 357452 16574 357480 149670
rect 360200 142860 360252 142866
rect 360200 142802 360252 142808
rect 360212 16574 360240 142802
rect 361578 18592 361634 18601
rect 361578 18527 361634 18536
rect 361592 16574 361620 18527
rect 374012 16574 374040 159287
rect 388536 158772 388588 158778
rect 388536 158714 388588 158720
rect 388548 158681 388576 158714
rect 376022 158672 376078 158681
rect 376022 158607 376024 158616
rect 376076 158607 376078 158616
rect 378598 158672 378654 158681
rect 378598 158607 378654 158616
rect 380990 158672 381046 158681
rect 380990 158607 381046 158616
rect 383566 158672 383622 158681
rect 383566 158607 383622 158616
rect 385958 158672 386014 158681
rect 385958 158607 386014 158616
rect 388534 158672 388590 158681
rect 388534 158607 388590 158616
rect 391478 158672 391534 158681
rect 391478 158607 391534 158616
rect 394238 158672 394294 158681
rect 394238 158607 394294 158616
rect 395894 158672 395950 158681
rect 395894 158607 395950 158616
rect 398470 158672 398526 158681
rect 398470 158607 398526 158616
rect 401046 158672 401102 158681
rect 401046 158607 401102 158616
rect 403990 158672 404046 158681
rect 403990 158607 404046 158616
rect 406474 158672 406530 158681
rect 406474 158607 406530 158616
rect 376024 158578 376076 158584
rect 378612 158574 378640 158607
rect 378600 158568 378652 158574
rect 378600 158510 378652 158516
rect 381004 158506 381032 158607
rect 380992 158500 381044 158506
rect 380992 158442 381044 158448
rect 383580 158438 383608 158607
rect 383568 158432 383620 158438
rect 383568 158374 383620 158380
rect 385972 158370 386000 158607
rect 385960 158364 386012 158370
rect 385960 158306 386012 158312
rect 391492 158302 391520 158607
rect 391480 158296 391532 158302
rect 391480 158238 391532 158244
rect 394252 158234 394280 158607
rect 394240 158228 394292 158234
rect 394240 158170 394292 158176
rect 395908 158166 395936 158607
rect 395896 158160 395948 158166
rect 395896 158102 395948 158108
rect 398484 158098 398512 158607
rect 398472 158092 398524 158098
rect 398472 158034 398524 158040
rect 401060 158030 401088 158607
rect 401048 158024 401100 158030
rect 401048 157966 401100 157972
rect 404004 157962 404032 158607
rect 403992 157956 404044 157962
rect 403992 157898 404044 157904
rect 406488 157894 406516 158607
rect 406476 157888 406528 157894
rect 406476 157830 406528 157836
rect 376760 152516 376812 152522
rect 376760 152458 376812 152464
rect 375378 80744 375434 80753
rect 375378 80679 375434 80688
rect 375392 16574 375420 80679
rect 376772 16574 376800 152458
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 357452 16546 357572 16574
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 374012 16546 374132 16574
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356336 4072 356388 4078
rect 356336 4014 356388 4020
rect 356348 480 356376 4014
rect 357544 480 357572 16546
rect 358728 6792 358780 6798
rect 358728 6734 358780 6740
rect 358740 480 358768 6734
rect 359924 4004 359976 4010
rect 359924 3946 359976 3952
rect 359936 480 359964 3946
rect 361132 480 361160 16546
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 372896 7608 372948 7614
rect 372896 7550 372948 7556
rect 369398 6896 369454 6905
rect 369398 6831 369454 6840
rect 367006 6624 367062 6633
rect 367006 6559 367062 6568
rect 365810 6080 365866 6089
rect 365810 6015 365866 6024
rect 364614 4992 364670 5001
rect 364614 4927 364670 4936
rect 363510 3224 363566 3233
rect 363510 3159 363566 3168
rect 363524 480 363552 3159
rect 364628 480 364656 4927
rect 365824 480 365852 6015
rect 367020 480 367048 6559
rect 368202 4856 368258 4865
rect 368202 4791 368258 4800
rect 368216 480 368244 4791
rect 369412 480 369440 6831
rect 370594 6488 370650 6497
rect 370594 6423 370650 6432
rect 370608 480 370636 6423
rect 371700 4140 371752 4146
rect 371700 4082 371752 4088
rect 371712 480 371740 4082
rect 372908 480 372936 7550
rect 374104 480 374132 16546
rect 375286 6760 375342 6769
rect 375286 6695 375342 6704
rect 375300 480 375328 6695
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 383566 9616 383622 9625
rect 383566 9551 383622 9560
rect 382372 6724 382424 6730
rect 382372 6666 382424 6672
rect 381176 3936 381228 3942
rect 379978 3904 380034 3913
rect 378876 3868 378928 3874
rect 381176 3878 381228 3884
rect 379978 3839 380034 3848
rect 378876 3810 378928 3816
rect 378888 480 378916 3810
rect 379992 480 380020 3839
rect 381188 480 381216 3878
rect 382384 480 382412 6666
rect 383580 480 383608 9551
rect 390650 9480 390706 9489
rect 390650 9415 390706 9424
rect 387154 8800 387210 8809
rect 387154 8735 387210 8744
rect 385960 6656 386012 6662
rect 385960 6598 386012 6604
rect 384762 4040 384818 4049
rect 384762 3975 384818 3984
rect 384776 480 384804 3975
rect 385972 480 386000 6598
rect 387168 480 387196 8735
rect 389454 6216 389510 6225
rect 389454 6151 389510 6160
rect 388260 3800 388312 3806
rect 388260 3742 388312 3748
rect 388272 480 388300 3742
rect 389468 480 389496 6151
rect 390664 480 390692 9415
rect 404818 9344 404874 9353
rect 404818 9279 404874 9288
rect 401324 8968 401376 8974
rect 401324 8910 401376 8916
rect 396540 6588 396592 6594
rect 396540 6530 396592 6536
rect 393042 6352 393098 6361
rect 393042 6287 393098 6296
rect 391846 3768 391902 3777
rect 391846 3703 391902 3712
rect 391860 480 391888 3703
rect 393056 480 393084 6287
rect 395344 3732 395396 3738
rect 395344 3674 395396 3680
rect 394238 3360 394294 3369
rect 394238 3295 394294 3304
rect 394252 480 394280 3295
rect 395356 480 395384 3674
rect 396552 480 396580 6530
rect 400128 6520 400180 6526
rect 400128 6462 400180 6468
rect 397734 3632 397790 3641
rect 397734 3567 397790 3576
rect 397748 480 397776 3567
rect 398930 3496 398986 3505
rect 398930 3431 398986 3440
rect 398944 480 398972 3431
rect 400140 480 400168 6462
rect 401336 480 401364 8910
rect 403624 6452 403676 6458
rect 403624 6394 403676 6400
rect 402520 3664 402572 3670
rect 402520 3606 402572 3612
rect 402532 480 402560 3606
rect 403636 480 403664 6394
rect 404832 480 404860 9279
rect 411902 9208 411958 9217
rect 411902 9143 411958 9152
rect 408406 9072 408462 9081
rect 408406 9007 408462 9016
rect 407212 6384 407264 6390
rect 407212 6326 407264 6332
rect 406016 3596 406068 3602
rect 406016 3538 406068 3544
rect 406028 480 406056 3538
rect 407224 480 407252 6326
rect 408420 480 408448 9007
rect 410800 6316 410852 6322
rect 410800 6258 410852 6264
rect 409604 3528 409656 3534
rect 409604 3470 409656 3476
rect 409616 480 409644 3470
rect 410812 480 410840 6258
rect 411916 480 411944 9143
rect 414294 8936 414350 8945
rect 414294 8871 414350 8880
rect 413100 3460 413152 3466
rect 413100 3402 413152 3408
rect 413112 480 413140 3402
rect 414308 480 414336 8871
rect 416688 6248 416740 6254
rect 416688 6190 416740 6196
rect 415492 3460 415544 3466
rect 415492 3402 415544 3408
rect 415504 480 415532 3402
rect 416700 480 416728 6190
rect 420184 6180 420236 6186
rect 420184 6122 420236 6128
rect 418988 3596 419040 3602
rect 418988 3538 419040 3544
rect 417884 3528 417936 3534
rect 417884 3470 417936 3476
rect 417896 480 417924 3470
rect 419000 480 419028 3538
rect 420196 480 420224 6122
rect 434444 4140 434496 4146
rect 434444 4082 434496 4088
rect 428464 4072 428516 4078
rect 428464 4014 428516 4020
rect 427268 4004 427320 4010
rect 427268 3946 427320 3952
rect 426164 3936 426216 3942
rect 426164 3878 426216 3884
rect 424968 3868 425020 3874
rect 424968 3810 425020 3816
rect 423772 3800 423824 3806
rect 423772 3742 423824 3748
rect 422576 3732 422628 3738
rect 422576 3674 422628 3680
rect 421380 3664 421432 3670
rect 421380 3606 421432 3612
rect 421392 480 421420 3606
rect 422588 480 422616 3674
rect 423784 480 423812 3742
rect 424980 480 425008 3810
rect 426176 480 426204 3878
rect 427280 480 427308 3946
rect 428476 480 428504 4014
rect 432050 3632 432106 3641
rect 432050 3567 432106 3576
rect 430856 3392 430908 3398
rect 429658 3360 429714 3369
rect 430856 3334 430908 3340
rect 429658 3295 429714 3304
rect 429672 480 429700 3295
rect 430868 480 430896 3334
rect 432064 480 432092 3567
rect 433248 3188 433300 3194
rect 433248 3130 433300 3136
rect 433260 480 433288 3130
rect 434456 480 434484 4082
rect 435548 3324 435600 3330
rect 435548 3266 435600 3272
rect 435560 480 435588 3266
rect 436756 480 436784 264386
rect 436848 158506 436876 308654
rect 436928 248328 436980 248334
rect 436928 248270 436980 248276
rect 436940 158778 436968 248270
rect 437480 248056 437532 248062
rect 437480 247998 437532 248004
rect 436928 158772 436980 158778
rect 436928 158714 436980 158720
rect 436836 158500 436888 158506
rect 436836 158442 436888 158448
rect 437492 3738 437520 247998
rect 437940 245608 437992 245614
rect 437940 245550 437992 245556
rect 437664 245540 437716 245546
rect 437664 245482 437716 245488
rect 437572 245268 437624 245274
rect 437572 245210 437624 245216
rect 437480 3732 437532 3738
rect 437480 3674 437532 3680
rect 437584 3466 437612 245210
rect 437676 3874 437704 245482
rect 437848 245404 437900 245410
rect 437848 245346 437900 245352
rect 437756 245200 437808 245206
rect 437756 245142 437808 245148
rect 437664 3868 437716 3874
rect 437664 3810 437716 3816
rect 437768 3534 437796 245142
rect 437860 3806 437888 245346
rect 437952 16574 437980 245550
rect 438044 158438 438072 308722
rect 439504 308644 439556 308650
rect 439504 308586 439556 308592
rect 438124 308508 438176 308514
rect 438124 308450 438176 308456
rect 438136 158642 438164 308450
rect 438216 248396 438268 248402
rect 438216 248338 438268 248344
rect 438124 158636 438176 158642
rect 438124 158578 438176 158584
rect 438032 158432 438084 158438
rect 438032 158374 438084 158380
rect 438228 157962 438256 248338
rect 438860 247988 438912 247994
rect 438860 247930 438912 247936
rect 438308 244860 438360 244866
rect 438308 244802 438360 244808
rect 438320 158302 438348 244802
rect 438308 158296 438360 158302
rect 438308 158238 438360 158244
rect 438216 157956 438268 157962
rect 438216 157898 438268 157904
rect 437952 16546 438072 16574
rect 437848 3800 437900 3806
rect 437848 3742 437900 3748
rect 437756 3528 437808 3534
rect 437756 3470 437808 3476
rect 437938 3496 437994 3505
rect 437572 3460 437624 3466
rect 437938 3431 437994 3440
rect 437572 3402 437624 3408
rect 437952 480 437980 3431
rect 438044 3398 438072 16546
rect 438872 3942 438900 247930
rect 439136 245472 439188 245478
rect 439136 245414 439188 245420
rect 438952 244996 439004 245002
rect 438952 244938 439004 244944
rect 438860 3936 438912 3942
rect 438860 3878 438912 3884
rect 438964 3602 438992 244938
rect 439044 244928 439096 244934
rect 439044 244870 439096 244876
rect 439056 3670 439084 244870
rect 439148 4146 439176 245414
rect 439320 245336 439372 245342
rect 439320 245278 439372 245284
rect 439228 245064 439280 245070
rect 439228 245006 439280 245012
rect 439136 4140 439188 4146
rect 439136 4082 439188 4088
rect 439240 4010 439268 245006
rect 439228 4004 439280 4010
rect 439228 3946 439280 3952
rect 439044 3664 439096 3670
rect 439044 3606 439096 3612
rect 438952 3596 439004 3602
rect 438952 3538 439004 3544
rect 439134 3496 439190 3505
rect 439134 3431 439190 3440
rect 438032 3392 438084 3398
rect 438032 3334 438084 3340
rect 439148 480 439176 3431
rect 439332 3330 439360 245278
rect 439412 245132 439464 245138
rect 439412 245074 439464 245080
rect 439424 4078 439452 245074
rect 439516 158370 439544 308586
rect 439596 308576 439648 308582
rect 439596 308518 439648 308524
rect 439608 158574 439636 308518
rect 440516 308440 440568 308446
rect 440516 308382 440568 308388
rect 440240 276752 440292 276758
rect 440240 276694 440292 276700
rect 439688 244792 439740 244798
rect 439688 244734 439740 244740
rect 439596 158568 439648 158574
rect 439596 158510 439648 158516
rect 439504 158364 439556 158370
rect 439504 158306 439556 158312
rect 439700 157894 439728 244734
rect 439688 157888 439740 157894
rect 439688 157830 439740 157836
rect 439412 4072 439464 4078
rect 439412 4014 439464 4020
rect 440252 3534 440280 276694
rect 440332 264376 440384 264382
rect 440332 264318 440384 264324
rect 440240 3528 440292 3534
rect 440240 3470 440292 3476
rect 439320 3324 439372 3330
rect 439320 3266 439372 3272
rect 440344 480 440372 264318
rect 440424 247920 440476 247926
rect 440424 247862 440476 247868
rect 440436 3194 440464 247862
rect 440528 158710 440556 308382
rect 445024 307216 445076 307222
rect 445024 307158 445076 307164
rect 442262 305960 442318 305969
rect 442262 305895 442318 305904
rect 441712 250776 441764 250782
rect 441712 250718 441764 250724
rect 441620 250708 441672 250714
rect 441620 250650 441672 250656
rect 440608 248192 440660 248198
rect 440608 248134 440660 248140
rect 440516 158704 440568 158710
rect 440516 158646 440568 158652
rect 440620 158234 440648 248134
rect 440608 158228 440660 158234
rect 440608 158170 440660 158176
rect 441632 16574 441660 250650
rect 441724 158098 441752 250718
rect 441804 248260 441856 248266
rect 441804 248202 441856 248208
rect 441712 158092 441764 158098
rect 441712 158034 441764 158040
rect 441816 158030 441844 248202
rect 441896 248124 441948 248130
rect 441896 248066 441948 248072
rect 441908 158166 441936 248066
rect 441896 158160 441948 158166
rect 441896 158102 441948 158108
rect 441804 158024 441856 158030
rect 441804 157966 441856 157972
rect 441632 16546 442212 16574
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 442184 3482 442212 16546
rect 442276 3670 442304 305895
rect 443644 304496 443696 304502
rect 443644 304438 443696 304444
rect 442264 3664 442316 3670
rect 442264 3606 442316 3612
rect 443656 3602 443684 304438
rect 444380 275460 444432 275466
rect 444380 275402 444432 275408
rect 444392 6914 444420 275402
rect 445036 16574 445064 307158
rect 445760 250640 445812 250646
rect 445760 250582 445812 250588
rect 445036 16546 445156 16574
rect 444392 6886 445064 6914
rect 443826 4040 443882 4049
rect 443826 3975 443882 3984
rect 443644 3596 443696 3602
rect 443644 3538 443696 3544
rect 440424 3188 440476 3194
rect 440424 3130 440476 3136
rect 441540 480 441568 3470
rect 442184 3454 442672 3482
rect 442644 480 442672 3454
rect 443840 480 443868 3975
rect 445036 480 445064 6886
rect 445128 3398 445156 16546
rect 445116 3392 445168 3398
rect 445116 3334 445168 3340
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 250582
rect 446416 73166 446444 443158
rect 458836 438190 458864 445810
rect 580356 445120 580408 445126
rect 580356 445062 580408 445068
rect 580264 445052 580316 445058
rect 580264 444994 580316 445000
rect 460204 444848 460256 444854
rect 460204 444790 460256 444796
rect 458824 438184 458876 438190
rect 458824 438126 458876 438132
rect 454040 298988 454092 298994
rect 454040 298930 454092 298936
rect 448520 287836 448572 287842
rect 448520 287778 448572 287784
rect 446404 73160 446456 73166
rect 446404 73102 446456 73108
rect 447416 3664 447468 3670
rect 447416 3606 447468 3612
rect 447428 480 447456 3606
rect 448532 3534 448560 287778
rect 449900 287768 449952 287774
rect 449900 287710 449952 287716
rect 448612 274168 448664 274174
rect 448612 274110 448664 274116
rect 448520 3528 448572 3534
rect 448520 3470 448572 3476
rect 448624 480 448652 274110
rect 449912 16574 449940 287710
rect 453304 284980 453356 284986
rect 453304 284922 453356 284928
rect 450544 271244 450596 271250
rect 450544 271186 450596 271192
rect 449912 16546 450492 16574
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 449820 480 449848 3470
rect 450464 3346 450492 16546
rect 450556 3466 450584 271186
rect 452660 258800 452712 258806
rect 452660 258742 452712 258748
rect 452672 16574 452700 258742
rect 452672 16546 453252 16574
rect 453224 3482 453252 16546
rect 453316 3602 453344 284922
rect 453304 3596 453356 3602
rect 453304 3538 453356 3544
rect 450544 3460 450596 3466
rect 450544 3402 450596 3408
rect 452108 3460 452160 3466
rect 453224 3454 453344 3482
rect 452108 3402 452160 3408
rect 450464 3318 450952 3346
rect 450924 480 450952 3318
rect 452120 480 452148 3402
rect 453316 480 453344 3454
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 298930
rect 456800 283756 456852 283762
rect 456800 283698 456852 283704
rect 456064 263016 456116 263022
rect 456064 262958 456116 262964
rect 456076 3670 456104 262958
rect 456064 3664 456116 3670
rect 456064 3606 456116 3612
rect 455696 3596 455748 3602
rect 455696 3538 455748 3544
rect 455708 480 455736 3538
rect 456812 3346 456840 283698
rect 459560 282260 459612 282266
rect 459560 282202 459612 282208
rect 458180 269952 458232 269958
rect 458180 269894 458232 269900
rect 456892 249212 456944 249218
rect 456892 249154 456944 249160
rect 456904 3466 456932 249154
rect 458192 16574 458220 269894
rect 459572 16574 459600 282202
rect 460216 113150 460244 444790
rect 494704 444780 494756 444786
rect 494704 444722 494756 444728
rect 462964 307148 463016 307154
rect 462964 307090 463016 307096
rect 462320 286544 462372 286550
rect 462320 286486 462372 286492
rect 460940 282328 460992 282334
rect 460940 282270 460992 282276
rect 460204 113144 460256 113150
rect 460204 113086 460256 113092
rect 460952 16574 460980 282270
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 456892 3460 456944 3466
rect 456892 3402 456944 3408
rect 458088 3460 458140 3466
rect 458088 3402 458140 3408
rect 456812 3318 456932 3346
rect 456904 480 456932 3318
rect 458100 480 458128 3402
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 286486
rect 462976 3738 463004 307090
rect 476762 305824 476818 305833
rect 476762 305759 476818 305768
rect 467104 296064 467156 296070
rect 467104 296006 467156 296012
rect 464344 268524 464396 268530
rect 464344 268466 464396 268472
rect 463700 264308 463752 264314
rect 463700 264250 463752 264256
rect 463712 16574 463740 264250
rect 463712 16546 464016 16574
rect 462964 3732 463016 3738
rect 462964 3674 463016 3680
rect 463988 480 464016 16546
rect 464356 3058 464384 268466
rect 466460 249144 466512 249150
rect 466460 249086 466512 249092
rect 466472 16574 466500 249086
rect 466472 16546 467052 16574
rect 465172 3664 465224 3670
rect 465172 3606 465224 3612
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 3606
rect 467024 3482 467052 16546
rect 467116 3602 467144 296006
rect 471244 294772 471296 294778
rect 471244 294714 471296 294720
rect 467840 286476 467892 286482
rect 467840 286418 467892 286424
rect 467852 16574 467880 286418
rect 467852 16546 468248 16574
rect 467104 3596 467156 3602
rect 467104 3538 467156 3544
rect 467024 3454 467512 3482
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 3454
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 469876 480 469904 3538
rect 471256 3534 471284 294714
rect 474740 280968 474792 280974
rect 474740 280910 474792 280916
rect 472624 280900 472676 280906
rect 472624 280842 472676 280848
rect 471980 254720 472032 254726
rect 471980 254662 472032 254668
rect 471992 16574 472020 254662
rect 471992 16546 472296 16574
rect 471060 3528 471112 3534
rect 471060 3470 471112 3476
rect 471244 3528 471296 3534
rect 471244 3470 471296 3476
rect 471072 480 471100 3470
rect 472268 480 472296 16546
rect 472636 3058 472664 280842
rect 474752 16574 474780 280910
rect 476120 267096 476172 267102
rect 476120 267038 476172 267044
rect 476132 16574 476160 267038
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 472624 3052 472676 3058
rect 472624 2994 472676 3000
rect 473464 480 473492 3470
rect 474556 3052 474608 3058
rect 474556 2994 474608 3000
rect 474568 480 474596 2994
rect 475764 480 475792 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 476776 3534 476804 305759
rect 485044 304428 485096 304434
rect 485044 304370 485096 304376
rect 481640 286408 481692 286414
rect 481640 286350 481692 286356
rect 477500 278180 477552 278186
rect 477500 278122 477552 278128
rect 477512 6914 477540 278122
rect 478144 254652 478196 254658
rect 478144 254594 478196 254600
rect 478156 16574 478184 254594
rect 478156 16546 478276 16574
rect 477512 6886 478184 6914
rect 476764 3528 476816 3534
rect 476764 3470 476816 3476
rect 478156 480 478184 6886
rect 478248 3262 478276 16546
rect 480536 3596 480588 3602
rect 480536 3538 480588 3544
rect 478236 3256 478288 3262
rect 478236 3198 478288 3204
rect 479340 3256 479392 3262
rect 479340 3198 479392 3204
rect 479352 480 479380 3198
rect 480548 480 480576 3538
rect 481652 3534 481680 286350
rect 481732 283688 481784 283694
rect 481732 283630 481784 283636
rect 481640 3528 481692 3534
rect 481640 3470 481692 3476
rect 481744 480 481772 283630
rect 484400 282192 484452 282198
rect 484400 282134 484452 282140
rect 484412 16574 484440 282134
rect 484412 16546 484808 16574
rect 484032 3596 484084 3602
rect 484032 3538 484084 3544
rect 482468 3528 482520 3534
rect 482468 3470 482520 3476
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3470
rect 484044 480 484072 3538
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 485056 3194 485084 304370
rect 489918 302832 489974 302841
rect 489918 302767 489974 302776
rect 485780 279540 485832 279546
rect 485780 279482 485832 279488
rect 485792 16574 485820 279482
rect 488540 265804 488592 265810
rect 488540 265746 488592 265752
rect 488552 16574 488580 265746
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 485044 3188 485096 3194
rect 485044 3130 485096 3136
rect 486436 480 486464 16546
rect 487620 3188 487672 3194
rect 487620 3130 487672 3136
rect 487632 480 487660 3130
rect 488828 480 488856 16546
rect 489932 3534 489960 302767
rect 491944 301640 491996 301646
rect 491944 301582 491996 301588
rect 491300 264240 491352 264246
rect 491300 264182 491352 264188
rect 490012 262948 490064 262954
rect 490012 262890 490064 262896
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 262890
rect 491312 16574 491340 264182
rect 491312 16546 491892 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 491864 3482 491892 16546
rect 491956 3602 491984 301582
rect 492680 261656 492732 261662
rect 492680 261598 492732 261604
rect 492692 16574 492720 261598
rect 494716 33114 494744 444722
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 500224 307080 500276 307086
rect 500224 307022 500276 307028
rect 498290 300112 498346 300121
rect 498290 300047 498346 300056
rect 496084 276684 496136 276690
rect 496084 276626 496136 276632
rect 495440 262880 495492 262886
rect 495440 262822 495492 262828
rect 494796 261588 494848 261594
rect 494796 261530 494848 261536
rect 494704 33108 494756 33114
rect 494704 33050 494756 33056
rect 492692 16546 493088 16574
rect 491944 3596 491996 3602
rect 491944 3538 491996 3544
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 491864 3454 492352 3482
rect 492324 480 492352 3454
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494704 3596 494756 3602
rect 494704 3538 494756 3544
rect 494716 480 494744 3538
rect 494808 2922 494836 261530
rect 494796 2916 494848 2922
rect 494796 2858 494848 2864
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 262822
rect 496096 3534 496124 276626
rect 498304 6914 498332 300047
rect 499580 275392 499632 275398
rect 499580 275334 499632 275340
rect 499592 16574 499620 275334
rect 499592 16546 500172 16574
rect 498212 6886 498332 6914
rect 496084 3528 496136 3534
rect 496084 3470 496136 3476
rect 497096 3528 497148 3534
rect 497096 3470 497148 3476
rect 497108 480 497136 3470
rect 498212 480 498240 6886
rect 500144 3482 500172 16546
rect 500236 3602 500264 307022
rect 511998 305688 512054 305697
rect 511998 305623 512054 305632
rect 502984 298920 503036 298926
rect 502984 298862 503036 298868
rect 502340 280832 502392 280838
rect 502340 280774 502392 280780
rect 502352 6914 502380 280774
rect 502996 16574 503024 298862
rect 507860 297560 507912 297566
rect 507860 297502 507912 297508
rect 506480 274100 506532 274106
rect 506480 274042 506532 274048
rect 503720 250572 503772 250578
rect 503720 250514 503772 250520
rect 502996 16546 503116 16574
rect 502352 6886 503024 6914
rect 500224 3596 500276 3602
rect 500224 3538 500276 3544
rect 501788 3596 501840 3602
rect 501788 3538 501840 3544
rect 500144 3454 500632 3482
rect 499396 2916 499448 2922
rect 499396 2858 499448 2864
rect 499408 480 499436 2858
rect 500604 480 500632 3454
rect 501800 480 501828 3538
rect 502996 480 503024 6886
rect 503088 3058 503116 16546
rect 503076 3052 503128 3058
rect 503076 2994 503128 3000
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 250514
rect 506492 3534 506520 274042
rect 506572 247852 506624 247858
rect 506572 247794 506624 247800
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506584 3346 506612 247794
rect 507872 16574 507900 297502
rect 511264 279472 511316 279478
rect 511264 279414 511316 279420
rect 509240 278112 509292 278118
rect 509240 278054 509292 278060
rect 509252 16574 509280 278054
rect 510620 252000 510672 252006
rect 510620 251942 510672 251948
rect 510632 16574 510660 251942
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511212 16574
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3318 506612 3346
rect 505376 3052 505428 3058
rect 505376 2994 505428 3000
rect 505388 480 505416 2994
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511184 3482 511212 16546
rect 511276 3602 511304 279414
rect 511264 3596 511316 3602
rect 511264 3538 511316 3544
rect 511184 3454 511304 3482
rect 511276 480 511304 3454
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 305623
rect 516784 304360 516836 304366
rect 516784 304302 516836 304308
rect 514024 295996 514076 296002
rect 514024 295938 514076 295944
rect 514036 3602 514064 295938
rect 514116 251932 514168 251938
rect 514116 251874 514168 251880
rect 513564 3596 513616 3602
rect 513564 3538 513616 3544
rect 514024 3596 514076 3602
rect 514024 3538 514076 3544
rect 513576 480 513604 3538
rect 514128 3534 514156 251874
rect 516138 245168 516194 245177
rect 516138 245103 516194 245112
rect 516152 16574 516180 245103
rect 516152 16546 516732 16574
rect 515956 3596 516008 3602
rect 515956 3538 516008 3544
rect 514116 3528 514168 3534
rect 514116 3470 514168 3476
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514772 480 514800 3470
rect 515968 480 515996 3538
rect 516704 3482 516732 16546
rect 516796 3874 516824 304302
rect 563704 304292 563756 304298
rect 563704 304234 563756 304240
rect 534724 301572 534776 301578
rect 534724 301514 534776 301520
rect 520280 298852 520332 298858
rect 520280 298794 520332 298800
rect 517520 247784 517572 247790
rect 517520 247726 517572 247732
rect 517532 16574 517560 247726
rect 517532 16546 517928 16574
rect 516784 3868 516836 3874
rect 516784 3810 516836 3816
rect 516704 3454 517192 3482
rect 517164 480 517192 3454
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 3868 519596 3874
rect 519544 3810 519596 3816
rect 519556 480 519584 3810
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 298794
rect 529940 294704 529992 294710
rect 529940 294646 529992 294652
rect 527824 293276 527876 293282
rect 527824 293218 527876 293224
rect 521660 272604 521712 272610
rect 521660 272546 521712 272552
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 272546
rect 527180 257440 527232 257446
rect 527180 257382 527232 257388
rect 523040 256012 523092 256018
rect 523040 255954 523092 255960
rect 523052 3534 523080 255954
rect 524420 246628 524472 246634
rect 524420 246570 524472 246576
rect 523130 245032 523186 245041
rect 523130 244967 523186 244976
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523144 3346 523172 244967
rect 524432 16574 524460 246570
rect 525800 246560 525852 246566
rect 525800 246502 525852 246508
rect 525812 16574 525840 246502
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523868 3528 523920 3534
rect 523868 3470 523920 3476
rect 523052 3318 523172 3346
rect 523052 480 523080 3318
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3470
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527192 6914 527220 257382
rect 527836 16574 527864 293218
rect 528560 269884 528612 269890
rect 528560 269826 528612 269832
rect 527836 16546 527956 16574
rect 527192 6886 527864 6914
rect 527836 480 527864 6886
rect 527928 3534 527956 16546
rect 527916 3528 527968 3534
rect 527916 3470 527968 3476
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 269826
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 294646
rect 531320 275324 531372 275330
rect 531320 275266 531372 275272
rect 531332 480 531360 275266
rect 534080 246492 534132 246498
rect 534080 246434 534132 246440
rect 531410 244896 531466 244905
rect 531410 244831 531466 244840
rect 531424 16574 531452 244831
rect 534092 16574 534120 246434
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3528 533764 3534
rect 533712 3470 533764 3476
rect 533724 480 533752 3470
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3194 534764 301514
rect 557540 298784 557592 298790
rect 557540 298726 557592 298732
rect 535460 294636 535512 294642
rect 535460 294578 535512 294584
rect 535472 6914 535500 294578
rect 538864 291848 538916 291854
rect 538864 291790 538916 291796
rect 536104 274032 536156 274038
rect 536104 273974 536156 273980
rect 536116 16574 536144 273974
rect 536116 16546 536236 16574
rect 535472 6886 536144 6914
rect 534724 3188 534776 3194
rect 534724 3130 534776 3136
rect 536116 480 536144 6886
rect 536208 4146 536236 16546
rect 536196 4140 536248 4146
rect 536196 4082 536248 4088
rect 538404 4140 538456 4146
rect 538404 4082 538456 4088
rect 537208 3188 537260 3194
rect 537208 3130 537260 3136
rect 537220 480 537248 3130
rect 538416 480 538444 4082
rect 538876 3058 538904 291790
rect 549904 290556 549956 290562
rect 549904 290498 549956 290504
rect 542360 278044 542412 278050
rect 542360 277986 542412 277992
rect 540244 271176 540296 271182
rect 540244 271118 540296 271124
rect 539692 268456 539744 268462
rect 539692 268398 539744 268404
rect 539704 6914 539732 268398
rect 539612 6886 539732 6914
rect 538864 3052 538916 3058
rect 538864 2994 538916 3000
rect 539612 480 539640 6886
rect 540256 2990 540284 271118
rect 542372 16574 542400 277986
rect 546500 261520 546552 261526
rect 546500 261462 546552 261468
rect 545120 250504 545172 250510
rect 545120 250446 545172 250452
rect 543740 246424 543792 246430
rect 543740 246366 543792 246372
rect 543752 16574 543780 246366
rect 545132 16574 545160 250446
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540796 3052 540848 3058
rect 540796 2994 540848 3000
rect 540244 2984 540296 2990
rect 540244 2926 540296 2932
rect 540808 480 540836 2994
rect 541992 2984 542044 2990
rect 541992 2926 542044 2932
rect 542004 480 542032 2926
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 261462
rect 549260 260160 549312 260166
rect 549260 260102 549312 260108
rect 547880 254584 547932 254590
rect 547880 254526 547932 254532
rect 547892 3534 547920 254526
rect 547972 247716 548024 247722
rect 547972 247658 548024 247664
rect 547880 3528 547932 3534
rect 547880 3470 547932 3476
rect 547984 3346 548012 247658
rect 549272 16574 549300 260102
rect 549272 16546 549852 16574
rect 548708 3528 548760 3534
rect 548708 3470 548760 3476
rect 549824 3482 549852 16546
rect 549916 3602 549944 290498
rect 552664 289196 552716 289202
rect 552664 289138 552716 289144
rect 552020 269816 552072 269822
rect 552020 269758 552072 269764
rect 552032 6914 552060 269758
rect 552676 16574 552704 289138
rect 556252 268388 556304 268394
rect 556252 268330 556304 268336
rect 554044 265736 554096 265742
rect 554044 265678 554096 265684
rect 553400 246356 553452 246362
rect 553400 246298 553452 246304
rect 553412 16574 553440 246298
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 552032 6886 552704 6914
rect 549904 3596 549956 3602
rect 549904 3538 549956 3544
rect 551468 3596 551520 3602
rect 551468 3538 551520 3544
rect 547892 3318 548012 3346
rect 547892 480 547920 3318
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 3470
rect 549824 3454 550312 3482
rect 550284 480 550312 3454
rect 551480 480 551508 3538
rect 552676 480 552704 6886
rect 552768 2990 552796 16546
rect 552756 2984 552808 2990
rect 552756 2926 552808 2932
rect 553780 480 553808 16546
rect 554056 3262 554084 265678
rect 556264 6914 556292 268330
rect 557552 16574 557580 298726
rect 560300 297492 560352 297498
rect 560300 297434 560352 297440
rect 558920 267028 558972 267034
rect 558920 266970 558972 266976
rect 558932 16574 558960 266970
rect 560312 16574 560340 297434
rect 561680 287700 561732 287706
rect 561680 287642 561732 287648
rect 560944 272536 560996 272542
rect 560944 272478 560996 272484
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 556172 6886 556292 6914
rect 554044 3256 554096 3262
rect 554044 3198 554096 3204
rect 554964 2984 555016 2990
rect 554964 2926 555016 2932
rect 554976 480 555004 2926
rect 556172 480 556200 6886
rect 557356 3256 557408 3262
rect 557356 3198 557408 3204
rect 557368 480 557396 3198
rect 558564 480 558592 16546
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 560956 3194 560984 272478
rect 561692 16574 561720 287642
rect 561692 16546 562088 16574
rect 560944 3188 560996 3194
rect 560944 3130 560996 3136
rect 562060 480 562088 16546
rect 563244 3188 563296 3194
rect 563244 3130 563296 3136
rect 563256 480 563284 3130
rect 563716 3058 563744 304234
rect 565820 301504 565872 301510
rect 565820 301446 565872 301452
rect 564532 251864 564584 251870
rect 564532 251806 564584 251812
rect 564544 6914 564572 251806
rect 565832 16574 565860 301446
rect 570604 297424 570656 297430
rect 570604 297366 570656 297372
rect 567200 290488 567252 290494
rect 567200 290430 567252 290436
rect 567212 16574 567240 290430
rect 567844 289128 567896 289134
rect 567844 289070 567896 289076
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 564452 6886 564572 6914
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 564452 480 564480 6886
rect 565636 3052 565688 3058
rect 565636 2994 565688 3000
rect 565648 480 565676 2994
rect 566844 480 566872 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3194 567884 289070
rect 570616 3466 570644 297366
rect 575480 286340 575532 286346
rect 575480 286282 575532 286288
rect 571340 283620 571392 283626
rect 571340 283562 571392 283568
rect 569132 3460 569184 3466
rect 569132 3402 569184 3408
rect 570604 3460 570656 3466
rect 570604 3402 570656 3408
rect 567844 3188 567896 3194
rect 567844 3130 567896 3136
rect 569144 480 569172 3402
rect 570328 3188 570380 3194
rect 570328 3130 570380 3136
rect 570340 480 570368 3130
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 283562
rect 574744 265668 574796 265674
rect 574744 265610 574796 265616
rect 574100 253292 574152 253298
rect 574100 253234 574152 253240
rect 571984 249076 572036 249082
rect 571984 249018 572036 249024
rect 571996 3534 572024 249018
rect 574112 16574 574140 253234
rect 574112 16546 574692 16574
rect 571984 3528 572036 3534
rect 571984 3470 572036 3476
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 574664 3482 574692 16546
rect 574756 3874 574784 265610
rect 575492 16574 575520 286282
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 578240 253224 578292 253230
rect 578240 253166 578292 253172
rect 578252 16574 578280 253166
rect 580276 152697 580304 444994
rect 580368 431633 580396 445062
rect 581000 439544 581052 439550
rect 581000 439486 581052 439492
rect 580354 431624 580410 431633
rect 580354 431559 580410 431568
rect 580448 260228 580500 260234
rect 580448 260170 580500 260176
rect 580356 258732 580408 258738
rect 580356 258674 580408 258680
rect 580368 192545 580396 258674
rect 580460 232393 580488 260170
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 574744 3868 574796 3874
rect 574744 3810 574796 3816
rect 572720 3460 572772 3466
rect 572720 3402 572772 3408
rect 572732 480 572760 3402
rect 573928 480 573956 3470
rect 574664 3454 575152 3482
rect 575124 480 575152 3454
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 3868 577464 3874
rect 577412 3810 577464 3816
rect 577424 480 577452 3810
rect 578620 480 578648 16546
rect 581012 3534 581040 439486
rect 582380 438184 582432 438190
rect 582380 438126 582432 438132
rect 581092 257372 581144 257378
rect 581092 257314 581144 257320
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581104 3346 581132 257314
rect 582392 16574 582420 438126
rect 582392 16546 583432 16574
rect 581828 3528 581880 3534
rect 581828 3470 581880 3476
rect 581012 3318 581132 3346
rect 581012 480 581040 3318
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581840 354 581868 3470
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581840 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3422 619112 3478 619168
rect 3330 579944 3386 580000
rect 3146 553832 3202 553888
rect 2962 527856 3018 527912
rect 2870 501744 2926 501800
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 2870 449520 2926 449576
rect 3514 606056 3570 606112
rect 3514 566888 3570 566944
rect 3606 514800 3662 514856
rect 217874 516840 217930 516896
rect 217782 515888 217838 515944
rect 217598 513712 217654 513768
rect 217322 488280 217378 488336
rect 217506 488008 217562 488064
rect 217690 489912 217746 489968
rect 3422 423580 3424 423600
rect 3424 423580 3476 423600
rect 3476 423580 3478 423600
rect 3422 423544 3478 423580
rect 2962 410488 3018 410544
rect 3330 397432 3386 397488
rect 3054 371320 3110 371376
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 2962 267144 3018 267200
rect 3146 254088 3202 254144
rect 3238 241032 3294 241088
rect 3330 214920 3386 214976
rect 3146 188808 3202 188864
rect 3146 110608 3202 110664
rect 3606 358400 3662 358456
rect 3514 201864 3570 201920
rect 3514 162832 3570 162888
rect 3606 149776 3662 149832
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3422 45464 3478 45520
rect 3422 6432 3478 6488
rect 219346 512760 219402 512816
rect 219254 510992 219310 511048
rect 219162 509904 219218 509960
rect 219070 508136 219126 508192
rect 242898 476856 242954 476912
rect 247038 476856 247094 476912
rect 238758 476740 238814 476776
rect 238758 476720 238760 476740
rect 238760 476720 238812 476740
rect 238812 476720 238814 476740
rect 97722 196832 97778 196888
rect 97814 195880 97870 195936
rect 97814 193704 97870 193760
rect 97538 192752 97594 192808
rect 97446 168272 97502 168328
rect 97630 190984 97686 191040
rect 97722 189896 97778 189952
rect 97906 188128 97962 188184
rect 97906 169904 97962 169960
rect 235998 476332 236054 476368
rect 235998 476312 236000 476332
rect 236000 476312 236052 476332
rect 236052 476312 236054 476332
rect 235998 476176 236054 476232
rect 237378 476196 237434 476232
rect 237378 476176 237380 476196
rect 237380 476176 237432 476196
rect 237432 476176 237434 476196
rect 240230 476176 240286 476232
rect 242806 476176 242862 476232
rect 244370 476448 244426 476504
rect 249798 477264 249854 477320
rect 268014 477264 268070 477320
rect 258078 476992 258134 477048
rect 252742 476856 252798 476912
rect 255410 476856 255466 476912
rect 244278 476332 244334 476368
rect 244278 476312 244280 476332
rect 244280 476312 244332 476332
rect 244332 476312 244334 476332
rect 245658 476196 245714 476232
rect 245658 476176 245660 476196
rect 245660 476176 245712 476196
rect 245712 476176 245714 476196
rect 247038 476176 247094 476232
rect 248510 476332 248566 476368
rect 248510 476312 248512 476332
rect 248512 476312 248564 476332
rect 248564 476312 248566 476332
rect 249890 476176 249946 476232
rect 252466 476312 252522 476368
rect 252650 476176 252706 476232
rect 253846 476196 253902 476232
rect 253846 476176 253848 476196
rect 253848 476176 253900 476196
rect 253900 476176 253902 476196
rect 255962 476312 256018 476368
rect 256606 476176 256662 476232
rect 258722 476720 258778 476776
rect 263598 476720 263654 476776
rect 258262 476584 258318 476640
rect 260838 476604 260894 476640
rect 260838 476584 260840 476604
rect 260840 476584 260892 476604
rect 260892 476584 260894 476604
rect 264242 476448 264298 476504
rect 264978 476448 265034 476504
rect 270498 476992 270554 477048
rect 304998 476992 305054 477048
rect 307758 476992 307814 477048
rect 261482 476312 261538 476368
rect 260746 476176 260802 476232
rect 262862 476176 262918 476232
rect 265622 476312 265678 476368
rect 267554 476312 267610 476368
rect 277950 476856 278006 476912
rect 302238 476856 302294 476912
rect 276018 476584 276074 476640
rect 266266 476176 266322 476232
rect 273258 476312 273314 476368
rect 274454 476312 274510 476368
rect 267646 476176 267702 476232
rect 269026 476176 269082 476232
rect 270406 476176 270462 476232
rect 271786 476176 271842 476232
rect 273166 476176 273222 476232
rect 274546 476176 274602 476232
rect 275926 476176 275982 476232
rect 277306 476176 277362 476232
rect 278686 476176 278742 476232
rect 280066 476176 280122 476232
rect 280250 476176 280306 476232
rect 283010 476176 283066 476232
rect 285770 476176 285826 476232
rect 287058 476176 287114 476232
rect 289910 476176 289966 476232
rect 292578 476176 292634 476232
rect 295430 476176 295486 476232
rect 298190 476176 298246 476232
rect 300950 476176 301006 476232
rect 310518 476856 310574 476912
rect 313278 476468 313334 476504
rect 313278 476448 313280 476468
rect 313280 476448 313332 476468
rect 313332 476448 313334 476468
rect 314658 476448 314714 476504
rect 322938 476856 322994 476912
rect 325790 476856 325846 476912
rect 317418 476332 317474 476368
rect 317418 476312 317420 476332
rect 317420 476312 317472 476332
rect 317472 476312 317474 476332
rect 320178 476312 320234 476368
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 484608 580226 484664
rect 238206 308352 238262 308408
rect 99286 168000 99342 168056
rect 153658 159840 153714 159896
rect 156050 159840 156106 159896
rect 160926 159840 160982 159896
rect 175922 159840 175978 159896
rect 165986 159568 166042 159624
rect 116214 158616 116270 158672
rect 118238 158616 118294 158672
rect 119894 158616 119950 158672
rect 120630 158616 120686 158672
rect 121918 158616 121974 158672
rect 126518 158636 126574 158672
rect 126518 158616 126520 158636
rect 126520 158616 126572 158636
rect 126572 158616 126574 158636
rect 117226 158072 117282 158128
rect 127622 158616 127678 158672
rect 200118 159296 200174 159352
rect 128726 158652 128728 158672
rect 128728 158652 128780 158672
rect 128780 158652 128782 158672
rect 128726 158616 128782 158652
rect 130566 158616 130622 158672
rect 131302 158616 131358 158672
rect 132406 158616 132462 158672
rect 133510 158616 133566 158672
rect 139306 158616 139362 158672
rect 159638 158616 159694 158672
rect 168286 158616 168342 158672
rect 188710 158616 188766 158672
rect 123942 158208 123998 158264
rect 135902 158480 135958 158536
rect 137006 158480 137062 158536
rect 138386 158480 138442 158536
rect 134614 158208 134670 158264
rect 124770 157528 124826 157584
rect 125414 157392 125470 157448
rect 133694 157392 133750 157448
rect 136086 157392 136142 157448
rect 133694 154400 133750 154456
rect 139674 158480 139730 158536
rect 141514 158208 141570 158264
rect 141790 158208 141846 158264
rect 146022 158208 146078 158264
rect 146390 158208 146446 158264
rect 150990 158208 151046 158264
rect 140686 157936 140742 157992
rect 139306 155896 139362 155952
rect 143078 157936 143134 157992
rect 144550 157936 144606 157992
rect 143998 157392 144054 157448
rect 145286 157664 145342 157720
rect 144550 155760 144606 155816
rect 136086 154264 136142 154320
rect 148690 158072 148746 158128
rect 148414 157664 148470 157720
rect 148782 157664 148838 157720
rect 149886 157392 149942 157448
rect 184018 158344 184074 158400
rect 185950 158344 186006 158400
rect 155774 157528 155830 157584
rect 151358 157392 151414 157448
rect 152646 157392 152702 157448
rect 153842 157392 153898 157448
rect 154486 157392 154542 157448
rect 151818 156576 151874 156632
rect 129738 153720 129794 153776
rect 157062 157392 157118 157448
rect 178038 156712 178094 156768
rect 160098 155216 160154 155272
rect 191470 158208 191526 158264
rect 195886 158208 195942 158264
rect 182178 155352 182234 155408
rect 198462 157392 198518 157448
rect 206006 158616 206062 158672
rect 201038 157528 201094 157584
rect 203430 157528 203486 157584
rect 207018 156848 207074 156904
rect 224958 155488 225014 155544
rect 238206 159160 238262 159216
rect 238298 158072 238354 158128
rect 241978 306312 242034 306368
rect 241978 306040 242034 306096
rect 250994 308624 251050 308680
rect 253386 155216 253442 155272
rect 254306 153720 254362 153776
rect 258446 156576 258502 156632
rect 260102 156712 260158 156768
rect 260102 141344 260158 141400
rect 262586 155352 262642 155408
rect 264334 148280 264390 148336
rect 265622 159296 265678 159352
rect 265162 128968 265218 129024
rect 268198 156848 268254 156904
rect 270498 306040 270554 306096
rect 270866 306040 270922 306096
rect 270958 155488 271014 155544
rect 272614 303048 272670 303104
rect 272614 155896 272670 155952
rect 272798 155760 272854 155816
rect 273902 147600 273958 147656
rect 276018 158344 276074 158400
rect 277490 307944 277546 308000
rect 277674 307808 277730 307864
rect 277122 158344 277178 158400
rect 276570 158072 276626 158128
rect 278778 307808 278834 307864
rect 279238 307808 279294 307864
rect 278686 300192 278742 300248
rect 278318 158208 278374 158264
rect 278686 158480 278742 158536
rect 279330 306176 279386 306232
rect 280066 306176 280122 306232
rect 279698 300600 279754 300656
rect 279790 300328 279846 300384
rect 281354 300464 281410 300520
rect 281078 157256 281134 157312
rect 283838 158208 283894 158264
rect 285494 307808 285550 307864
rect 285126 157528 285182 157584
rect 286782 247016 286838 247072
rect 287886 247016 287942 247072
rect 288070 247016 288126 247072
rect 288990 247016 289046 247072
rect 289174 247016 289230 247072
rect 289266 158752 289322 158808
rect 289450 155760 289506 155816
rect 289358 153040 289414 153096
rect 289634 155896 289690 155952
rect 290646 247016 290702 247072
rect 290738 156576 290794 156632
rect 291014 245112 291070 245168
rect 290922 157936 290978 157992
rect 290922 156712 290978 156768
rect 291750 244332 291752 244352
rect 291752 244332 291804 244352
rect 291804 244332 291806 244352
rect 291750 244296 291806 244332
rect 292210 244296 292266 244352
rect 292118 196016 292174 196072
rect 292394 247016 292450 247072
rect 292394 166232 292450 166288
rect 293406 244432 293462 244488
rect 293498 158752 293554 158808
rect 293682 244296 293738 244352
rect 293866 158888 293922 158944
rect 295062 157392 295118 157448
rect 295246 244704 295302 244760
rect 296626 307808 296682 307864
rect 296994 308216 297050 308272
rect 297270 307944 297326 308000
rect 298098 309032 298154 309088
rect 297914 308080 297970 308136
rect 297638 307808 297694 307864
rect 296810 246200 296866 246256
rect 296718 244840 296774 244896
rect 297270 195880 297326 195936
rect 297362 192752 297418 192808
rect 297270 191664 297326 191720
rect 297270 190984 297326 191040
rect 297086 189896 297142 189952
rect 297086 189080 297142 189136
rect 297178 169904 297234 169960
rect 297454 191664 297510 191720
rect 297454 189080 297510 189136
rect 297730 168272 297786 168328
rect 297638 168000 297694 168056
rect 299202 307944 299258 308000
rect 299018 307808 299074 307864
rect 298374 244296 298430 244352
rect 298742 244296 298798 244352
rect 298282 159296 298338 159352
rect 299294 245520 299350 245576
rect 298742 188128 298798 188184
rect 298926 196832 298982 196888
rect 299110 193704 299166 193760
rect 299110 187720 299166 187776
rect 299018 158752 299074 158808
rect 299846 248104 299902 248160
rect 299938 247968 299994 248024
rect 300674 247968 300730 248024
rect 299754 244568 299810 244624
rect 300950 245248 301006 245304
rect 301226 247560 301282 247616
rect 301318 247288 301374 247344
rect 302330 245384 302386 245440
rect 302422 245112 302478 245168
rect 302606 247696 302662 247752
rect 302790 247832 302846 247888
rect 302698 247424 302754 247480
rect 305274 247968 305330 248024
rect 302514 244976 302570 245032
rect 306562 245520 306618 245576
rect 308126 247560 308182 247616
rect 311622 302912 311678 302968
rect 310978 298696 311034 298752
rect 310886 287680 310942 287736
rect 312634 305904 312690 305960
rect 316130 307808 316186 307864
rect 318154 307808 318210 307864
rect 318982 306312 319038 306368
rect 320086 306312 320142 306368
rect 320086 305768 320142 305824
rect 321098 302776 321154 302832
rect 321926 300056 321982 300112
rect 324226 305632 324282 305688
rect 309230 245248 309286 245304
rect 324410 305496 324466 305552
rect 324594 305496 324650 305552
rect 324318 245112 324374 245168
rect 325698 244976 325754 245032
rect 331402 305496 331458 305552
rect 331678 305496 331734 305552
rect 327078 244840 327134 244896
rect 301042 244704 301098 244760
rect 337934 308352 337990 308408
rect 338946 306176 339002 306232
rect 340050 303320 340106 303376
rect 341062 303184 341118 303240
rect 342442 303048 342498 303104
rect 347042 308624 347098 308680
rect 348330 308896 348386 308952
rect 349618 308760 349674 308816
rect 352286 308488 352342 308544
rect 353390 306040 353446 306096
rect 352654 300600 352710 300656
rect 355782 300328 355838 300384
rect 356426 300464 356482 300520
rect 359186 300192 359242 300248
rect 348238 159840 348294 159896
rect 350998 159840 351054 159896
rect 356058 159840 356114 159896
rect 358450 159840 358506 159896
rect 360934 159840 360990 159896
rect 368294 159840 368350 159896
rect 300858 152360 300914 152416
rect 316038 158616 316094 158672
rect 317050 158616 317106 158672
rect 319442 158616 319498 158672
rect 320546 158616 320602 158672
rect 321650 158616 321706 158672
rect 323122 158616 323178 158672
rect 324226 157800 324282 157856
rect 324870 157392 324926 157448
rect 327538 158616 327594 158672
rect 328274 158616 328330 158672
rect 329930 158616 329986 158672
rect 330298 158616 330354 158672
rect 331218 158636 331274 158672
rect 331218 158616 331220 158636
rect 331220 158616 331272 158636
rect 331272 158616 331274 158636
rect 332322 158616 332378 158672
rect 333610 158616 333666 158672
rect 334530 158616 334586 158672
rect 335818 158616 335874 158672
rect 336002 158616 336058 158672
rect 336922 158616 336978 158672
rect 338394 158652 338396 158672
rect 338396 158652 338448 158672
rect 338448 158652 338450 158672
rect 338394 158616 338450 158652
rect 338118 158208 338174 158264
rect 353574 159568 353630 159624
rect 365902 159568 365958 159624
rect 373998 159296 374054 159352
rect 339314 158616 339370 158672
rect 340970 158616 341026 158672
rect 343546 158616 343602 158672
rect 347594 158616 347650 158672
rect 354402 158616 354458 158672
rect 355230 158616 355286 158672
rect 356978 158616 357034 158672
rect 363418 158616 363474 158672
rect 370962 158616 371018 158672
rect 373446 158652 373448 158672
rect 373448 158652 373500 158672
rect 373500 158652 373502 158672
rect 373446 158616 373502 158652
rect 343914 158208 343970 158264
rect 341154 157936 341210 157992
rect 339590 157800 339646 157856
rect 342350 157800 342406 157856
rect 345110 157936 345166 157992
rect 346398 157936 346454 157992
rect 345754 157392 345810 157448
rect 348698 158208 348754 158264
rect 353298 158208 353354 158264
rect 349802 157392 349858 157448
rect 351090 157392 351146 157448
rect 352194 157392 352250 157448
rect 361578 18536 361634 18592
rect 376022 158636 376078 158672
rect 376022 158616 376024 158636
rect 376024 158616 376076 158636
rect 376076 158616 376078 158636
rect 378598 158616 378654 158672
rect 380990 158616 381046 158672
rect 383566 158616 383622 158672
rect 385958 158616 386014 158672
rect 388534 158616 388590 158672
rect 391478 158616 391534 158672
rect 394238 158616 394294 158672
rect 395894 158616 395950 158672
rect 398470 158616 398526 158672
rect 401046 158616 401102 158672
rect 403990 158616 404046 158672
rect 406474 158616 406530 158672
rect 375378 80688 375434 80744
rect 369398 6840 369454 6896
rect 367006 6568 367062 6624
rect 365810 6024 365866 6080
rect 364614 4936 364670 4992
rect 363510 3168 363566 3224
rect 368202 4800 368258 4856
rect 370594 6432 370650 6488
rect 375286 6704 375342 6760
rect 383566 9560 383622 9616
rect 379978 3848 380034 3904
rect 390650 9424 390706 9480
rect 387154 8744 387210 8800
rect 384762 3984 384818 4040
rect 389454 6160 389510 6216
rect 404818 9288 404874 9344
rect 393042 6296 393098 6352
rect 391846 3712 391902 3768
rect 394238 3304 394294 3360
rect 397734 3576 397790 3632
rect 398930 3440 398986 3496
rect 411902 9152 411958 9208
rect 408406 9016 408462 9072
rect 414294 8880 414350 8936
rect 432050 3576 432106 3632
rect 429658 3304 429714 3360
rect 437938 3440 437994 3496
rect 439134 3440 439190 3496
rect 442262 305904 442318 305960
rect 443826 3984 443882 4040
rect 476762 305768 476818 305824
rect 489918 302776 489974 302832
rect 580170 378392 580226 378448
rect 579894 325216 579950 325272
rect 498290 300056 498346 300112
rect 511998 305632 512054 305688
rect 516138 245112 516194 245168
rect 523130 244976 523186 245032
rect 531410 244840 531466 244896
rect 579894 272176 579950 272232
rect 580354 431568 580410 431624
rect 580446 232328 580502 232384
rect 580354 192480 580410 192536
rect 580262 152632 580318 152688
rect 579802 112784 579858 112840
rect 580170 72936 580226 72992
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 583520 524364 584960 524604
rect 217869 516898 217935 516901
rect 219390 516898 220064 516924
rect 217869 516896 220064 516898
rect 217869 516840 217874 516896
rect 217930 516864 220064 516896
rect 217930 516840 219450 516864
rect 217869 516838 219450 516840
rect 217869 516835 217935 516838
rect 217777 515946 217843 515949
rect 219390 515946 220064 515972
rect 217777 515944 220064 515946
rect 217777 515888 217782 515944
rect 217838 515912 220064 515944
rect 217838 515888 219450 515912
rect 217777 515886 219450 515888
rect 217777 515883 217843 515886
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 217593 513770 217659 513773
rect 219390 513770 220064 513796
rect 217593 513768 220064 513770
rect 217593 513712 217598 513768
rect 217654 513736 220064 513768
rect 217654 513712 219450 513736
rect 217593 513710 219450 513712
rect 217593 513707 217659 513710
rect 219390 512821 220064 512844
rect 219341 512816 220064 512821
rect 219341 512760 219346 512816
rect 219402 512784 220064 512816
rect 219402 512760 219450 512784
rect 219341 512758 219450 512760
rect 219341 512755 219407 512758
rect 583520 511172 584960 511412
rect 219249 511050 219315 511053
rect 219390 511050 220064 511076
rect 219249 511048 220064 511050
rect 219249 510992 219254 511048
rect 219310 511016 220064 511048
rect 219310 510992 219450 511016
rect 219249 510990 219450 510992
rect 219249 510987 219315 510990
rect 219157 509962 219223 509965
rect 219390 509962 220064 509988
rect 219157 509960 220064 509962
rect 219157 509904 219162 509960
rect 219218 509928 220064 509960
rect 219218 509904 219450 509928
rect 219157 509902 219450 509904
rect 219157 509899 219223 509902
rect 219065 508194 219131 508197
rect 219390 508194 220064 508220
rect 219065 508192 220064 508194
rect 219065 508136 219070 508192
rect 219126 508160 220064 508192
rect 219126 508136 219450 508160
rect 219065 508134 219450 508136
rect 219065 508131 219131 508134
rect -960 501802 480 501892
rect 2865 501802 2931 501805
rect -960 501800 2931 501802
rect -960 501744 2870 501800
rect 2926 501744 2931 501800
rect -960 501742 2931 501744
rect -960 501652 480 501742
rect 2865 501739 2931 501742
rect 583520 497844 584960 498084
rect 217685 489970 217751 489973
rect 219390 489970 220064 489996
rect 217685 489968 220064 489970
rect 217685 489912 217690 489968
rect 217746 489936 220064 489968
rect 217746 489912 219450 489936
rect 217685 489910 219450 489912
rect 217685 489907 217751 489910
rect -960 488596 480 488836
rect 217317 488338 217383 488341
rect 219390 488338 220064 488364
rect 217317 488336 220064 488338
rect 217317 488280 217322 488336
rect 217378 488304 220064 488336
rect 217378 488280 219450 488304
rect 217317 488278 219450 488280
rect 217317 488275 217383 488278
rect 217501 488066 217567 488069
rect 219390 488066 220064 488092
rect 217501 488064 220064 488066
rect 217501 488008 217506 488064
rect 217562 488032 220064 488064
rect 217562 488008 219450 488032
rect 217501 488006 219450 488008
rect 217501 488003 217567 488006
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 249793 477322 249859 477325
rect 250662 477322 250668 477324
rect 249793 477320 250668 477322
rect 249793 477264 249798 477320
rect 249854 477264 250668 477320
rect 249793 477262 250668 477264
rect 249793 477259 249859 477262
rect 250662 477260 250668 477262
rect 250732 477260 250738 477324
rect 268009 477322 268075 477325
rect 268326 477322 268332 477324
rect 268009 477320 268332 477322
rect 268009 477264 268014 477320
rect 268070 477264 268332 477320
rect 268009 477262 268332 477264
rect 268009 477259 268075 477262
rect 268326 477260 268332 477262
rect 268396 477260 268402 477324
rect 258073 477052 258139 477053
rect 258022 476988 258028 477052
rect 258092 477050 258139 477052
rect 270493 477050 270559 477053
rect 270902 477050 270908 477052
rect 258092 477048 258184 477050
rect 258134 476992 258184 477048
rect 258092 476990 258184 476992
rect 270493 477048 270908 477050
rect 270493 476992 270498 477048
rect 270554 476992 270908 477048
rect 270493 476990 270908 476992
rect 258092 476988 258139 476990
rect 258073 476987 258139 476988
rect 270493 476987 270559 476990
rect 270902 476988 270908 476990
rect 270972 476988 270978 477052
rect 304993 477050 305059 477053
rect 305862 477050 305868 477052
rect 304993 477048 305868 477050
rect 304993 476992 304998 477048
rect 305054 476992 305868 477048
rect 304993 476990 305868 476992
rect 304993 476987 305059 476990
rect 305862 476988 305868 476990
rect 305932 476988 305938 477052
rect 307753 477050 307819 477053
rect 308438 477050 308444 477052
rect 307753 477048 308444 477050
rect 307753 476992 307758 477048
rect 307814 476992 308444 477048
rect 307753 476990 308444 476992
rect 307753 476987 307819 476990
rect 308438 476988 308444 476990
rect 308508 476988 308514 477052
rect 242893 476914 242959 476917
rect 243118 476914 243124 476916
rect 242893 476912 243124 476914
rect 242893 476856 242898 476912
rect 242954 476856 243124 476912
rect 242893 476854 243124 476856
rect 242893 476851 242959 476854
rect 243118 476852 243124 476854
rect 243188 476852 243194 476916
rect 247033 476914 247099 476917
rect 248270 476914 248276 476916
rect 247033 476912 248276 476914
rect 247033 476856 247038 476912
rect 247094 476856 248276 476912
rect 247033 476854 248276 476856
rect 247033 476851 247099 476854
rect 248270 476852 248276 476854
rect 248340 476852 248346 476916
rect 252737 476914 252803 476917
rect 253606 476914 253612 476916
rect 252737 476912 253612 476914
rect 252737 476856 252742 476912
rect 252798 476856 253612 476912
rect 252737 476854 253612 476856
rect 252737 476851 252803 476854
rect 253606 476852 253612 476854
rect 253676 476852 253682 476916
rect 255405 476914 255471 476917
rect 256182 476914 256188 476916
rect 255405 476912 256188 476914
rect 255405 476856 255410 476912
rect 255466 476856 256188 476912
rect 255405 476854 256188 476856
rect 255405 476851 255471 476854
rect 256182 476852 256188 476854
rect 256252 476852 256258 476916
rect 277945 476914 278011 476917
rect 278446 476914 278452 476916
rect 277945 476912 278452 476914
rect 277945 476856 277950 476912
rect 278006 476856 278452 476912
rect 277945 476854 278452 476856
rect 277945 476851 278011 476854
rect 278446 476852 278452 476854
rect 278516 476852 278522 476916
rect 302233 476914 302299 476917
rect 303470 476914 303476 476916
rect 302233 476912 303476 476914
rect 302233 476856 302238 476912
rect 302294 476856 303476 476912
rect 302233 476854 303476 476856
rect 302233 476851 302299 476854
rect 303470 476852 303476 476854
rect 303540 476852 303546 476916
rect 310513 476914 310579 476917
rect 311014 476914 311020 476916
rect 310513 476912 311020 476914
rect 310513 476856 310518 476912
rect 310574 476856 311020 476912
rect 310513 476854 311020 476856
rect 310513 476851 310579 476854
rect 311014 476852 311020 476854
rect 311084 476852 311090 476916
rect 322933 476914 322999 476917
rect 323342 476914 323348 476916
rect 322933 476912 323348 476914
rect 322933 476856 322938 476912
rect 322994 476856 323348 476912
rect 322933 476854 323348 476856
rect 322933 476851 322999 476854
rect 323342 476852 323348 476854
rect 323412 476852 323418 476916
rect 325785 476914 325851 476917
rect 325918 476914 325924 476916
rect 325785 476912 325924 476914
rect 325785 476856 325790 476912
rect 325846 476856 325924 476912
rect 325785 476854 325924 476856
rect 325785 476851 325851 476854
rect 325918 476852 325924 476854
rect 325988 476852 325994 476916
rect 238753 476778 238819 476781
rect 239622 476778 239628 476780
rect 238753 476776 239628 476778
rect 238753 476720 238758 476776
rect 238814 476720 239628 476776
rect 238753 476718 239628 476720
rect 238753 476715 238819 476718
rect 239622 476716 239628 476718
rect 239692 476716 239698 476780
rect 257102 476716 257108 476780
rect 257172 476778 257178 476780
rect 258717 476778 258783 476781
rect 263593 476780 263659 476781
rect 257172 476776 258783 476778
rect 257172 476720 258722 476776
rect 258778 476720 258783 476776
rect 257172 476718 258783 476720
rect 257172 476716 257178 476718
rect 258717 476715 258783 476718
rect 263542 476716 263548 476780
rect 263612 476778 263659 476780
rect 263612 476776 263704 476778
rect 263654 476720 263704 476776
rect 263612 476718 263704 476720
rect 263612 476716 263659 476718
rect 263593 476715 263659 476716
rect 258257 476642 258323 476645
rect 258390 476642 258396 476644
rect 258257 476640 258396 476642
rect 258257 476584 258262 476640
rect 258318 476584 258396 476640
rect 258257 476582 258396 476584
rect 258257 476579 258323 476582
rect 258390 476580 258396 476582
rect 258460 476580 258466 476644
rect 260833 476642 260899 476645
rect 276013 476644 276079 476645
rect 260966 476642 260972 476644
rect 260833 476640 260972 476642
rect 260833 476584 260838 476640
rect 260894 476584 260972 476640
rect 260833 476582 260972 476584
rect 260833 476579 260899 476582
rect 260966 476580 260972 476582
rect 261036 476580 261042 476644
rect 276013 476642 276060 476644
rect 275968 476640 276060 476642
rect 275968 476584 276018 476640
rect 275968 476582 276060 476584
rect 276013 476580 276060 476582
rect 276124 476580 276130 476644
rect 276013 476579 276079 476580
rect 244365 476506 244431 476509
rect 245326 476506 245332 476508
rect 244365 476504 245332 476506
rect 244365 476448 244370 476504
rect 244426 476448 245332 476504
rect 244365 476446 245332 476448
rect 244365 476443 244431 476446
rect 245326 476444 245332 476446
rect 245396 476444 245402 476508
rect 262806 476444 262812 476508
rect 262876 476506 262882 476508
rect 264237 476506 264303 476509
rect 262876 476504 264303 476506
rect 262876 476448 264242 476504
rect 264298 476448 264303 476504
rect 262876 476446 264303 476448
rect 262876 476444 262882 476446
rect 264237 476443 264303 476446
rect 264973 476506 265039 476509
rect 265934 476506 265940 476508
rect 264973 476504 265940 476506
rect 264973 476448 264978 476504
rect 265034 476448 265940 476504
rect 264973 476446 265940 476448
rect 264973 476443 265039 476446
rect 265934 476444 265940 476446
rect 266004 476444 266010 476508
rect 313273 476506 313339 476509
rect 313406 476506 313412 476508
rect 313273 476504 313412 476506
rect 313273 476448 313278 476504
rect 313334 476448 313412 476504
rect 313273 476446 313412 476448
rect 313273 476443 313339 476446
rect 313406 476444 313412 476446
rect 313476 476444 313482 476508
rect 314653 476506 314719 476509
rect 315798 476506 315804 476508
rect 314653 476504 315804 476506
rect 314653 476448 314658 476504
rect 314714 476448 315804 476504
rect 314653 476446 315804 476448
rect 314653 476443 314719 476446
rect 315798 476444 315804 476446
rect 315868 476444 315874 476508
rect 235993 476372 236059 476373
rect 244273 476372 244339 476373
rect 235942 476308 235948 476372
rect 236012 476370 236059 476372
rect 236012 476368 236104 476370
rect 236054 476312 236104 476368
rect 236012 476310 236104 476312
rect 236012 476308 236059 476310
rect 244222 476308 244228 476372
rect 244292 476370 244339 476372
rect 248505 476370 248571 476373
rect 248638 476370 248644 476372
rect 244292 476368 244384 476370
rect 244334 476312 244384 476368
rect 244292 476310 244384 476312
rect 248505 476368 248644 476370
rect 248505 476312 248510 476368
rect 248566 476312 248644 476368
rect 248505 476310 248644 476312
rect 244292 476308 244339 476310
rect 235993 476307 236059 476308
rect 244273 476307 244339 476308
rect 248505 476307 248571 476310
rect 248638 476308 248644 476310
rect 248708 476308 248714 476372
rect 252318 476308 252324 476372
rect 252388 476370 252394 476372
rect 252461 476370 252527 476373
rect 252388 476368 252527 476370
rect 252388 476312 252466 476368
rect 252522 476312 252527 476368
rect 252388 476310 252527 476312
rect 252388 476308 252394 476310
rect 252461 476307 252527 476310
rect 254526 476308 254532 476372
rect 254596 476370 254602 476372
rect 255957 476370 256023 476373
rect 254596 476368 256023 476370
rect 254596 476312 255962 476368
rect 256018 476312 256023 476368
rect 254596 476310 256023 476312
rect 254596 476308 254602 476310
rect 255957 476307 256023 476310
rect 260782 476308 260788 476372
rect 260852 476370 260858 476372
rect 261477 476370 261543 476373
rect 260852 476368 261543 476370
rect 260852 476312 261482 476368
rect 261538 476312 261543 476368
rect 260852 476310 261543 476312
rect 260852 476308 260858 476310
rect 261477 476307 261543 476310
rect 263910 476308 263916 476372
rect 263980 476370 263986 476372
rect 265617 476370 265683 476373
rect 267549 476372 267615 476373
rect 267549 476370 267596 476372
rect 263980 476368 265683 476370
rect 263980 476312 265622 476368
rect 265678 476312 265683 476368
rect 263980 476310 265683 476312
rect 267504 476368 267596 476370
rect 267504 476312 267554 476368
rect 267504 476310 267596 476312
rect 263980 476308 263986 476310
rect 265617 476307 265683 476310
rect 267549 476308 267596 476310
rect 267660 476308 267666 476372
rect 273253 476370 273319 476373
rect 274449 476372 274515 476373
rect 273478 476370 273484 476372
rect 273253 476368 273484 476370
rect 273253 476312 273258 476368
rect 273314 476312 273484 476368
rect 273253 476310 273484 476312
rect 267549 476307 267615 476308
rect 273253 476307 273319 476310
rect 273478 476308 273484 476310
rect 273548 476308 273554 476372
rect 274398 476308 274404 476372
rect 274468 476370 274515 476372
rect 317413 476370 317479 476373
rect 318374 476370 318380 476372
rect 274468 476368 274560 476370
rect 274510 476312 274560 476368
rect 274468 476310 274560 476312
rect 317413 476368 318380 476370
rect 317413 476312 317418 476368
rect 317474 476312 318380 476368
rect 317413 476310 318380 476312
rect 274468 476308 274515 476310
rect 274449 476307 274515 476308
rect 317413 476307 317479 476310
rect 318374 476308 318380 476310
rect 318444 476308 318450 476372
rect 320173 476370 320239 476373
rect 320950 476370 320956 476372
rect 320173 476368 320956 476370
rect 320173 476312 320178 476368
rect 320234 476312 320956 476368
rect 320173 476310 320956 476312
rect 320173 476307 320239 476310
rect 320950 476308 320956 476310
rect 321020 476308 321026 476372
rect 235993 476234 236059 476237
rect 237046 476234 237052 476236
rect 235993 476232 237052 476234
rect 235993 476176 235998 476232
rect 236054 476176 237052 476232
rect 235993 476174 237052 476176
rect 235993 476171 236059 476174
rect 237046 476172 237052 476174
rect 237116 476172 237122 476236
rect 237373 476234 237439 476237
rect 238150 476234 238156 476236
rect 237373 476232 238156 476234
rect 237373 476176 237378 476232
rect 237434 476176 238156 476232
rect 237373 476174 238156 476176
rect 237373 476171 237439 476174
rect 238150 476172 238156 476174
rect 238220 476172 238226 476236
rect 240225 476234 240291 476237
rect 240542 476234 240548 476236
rect 240225 476232 240548 476234
rect 240225 476176 240230 476232
rect 240286 476176 240548 476232
rect 240225 476174 240548 476176
rect 240225 476171 240291 476174
rect 240542 476172 240548 476174
rect 240612 476172 240618 476236
rect 241830 476172 241836 476236
rect 241900 476234 241906 476236
rect 242801 476234 242867 476237
rect 241900 476232 242867 476234
rect 241900 476176 242806 476232
rect 242862 476176 242867 476232
rect 241900 476174 242867 476176
rect 241900 476172 241906 476174
rect 242801 476171 242867 476174
rect 245653 476234 245719 476237
rect 246430 476234 246436 476236
rect 245653 476232 246436 476234
rect 245653 476176 245658 476232
rect 245714 476176 246436 476232
rect 245653 476174 246436 476176
rect 245653 476171 245719 476174
rect 246430 476172 246436 476174
rect 246500 476172 246506 476236
rect 247033 476234 247099 476237
rect 247534 476234 247540 476236
rect 247033 476232 247540 476234
rect 247033 476176 247038 476232
rect 247094 476176 247540 476232
rect 247033 476174 247540 476176
rect 247033 476171 247099 476174
rect 247534 476172 247540 476174
rect 247604 476172 247610 476236
rect 249885 476234 249951 476237
rect 250110 476234 250116 476236
rect 249885 476232 250116 476234
rect 249885 476176 249890 476232
rect 249946 476176 250116 476232
rect 249885 476174 250116 476176
rect 249885 476171 249951 476174
rect 250110 476172 250116 476174
rect 250180 476172 250186 476236
rect 251398 476172 251404 476236
rect 251468 476234 251474 476236
rect 252645 476234 252711 476237
rect 251468 476232 252711 476234
rect 251468 476176 252650 476232
rect 252706 476176 252711 476232
rect 251468 476174 252711 476176
rect 251468 476172 251474 476174
rect 252645 476171 252711 476174
rect 253422 476172 253428 476236
rect 253492 476234 253498 476236
rect 253841 476234 253907 476237
rect 253492 476232 253907 476234
rect 253492 476176 253846 476232
rect 253902 476176 253907 476232
rect 253492 476174 253907 476176
rect 253492 476172 253498 476174
rect 253841 476171 253907 476174
rect 255814 476172 255820 476236
rect 255884 476234 255890 476236
rect 256601 476234 256667 476237
rect 255884 476232 256667 476234
rect 255884 476176 256606 476232
rect 256662 476176 256667 476232
rect 255884 476174 256667 476176
rect 255884 476172 255890 476174
rect 256601 476171 256667 476174
rect 259494 476172 259500 476236
rect 259564 476234 259570 476236
rect 260741 476234 260807 476237
rect 259564 476232 260807 476234
rect 259564 476176 260746 476232
rect 260802 476176 260807 476232
rect 259564 476174 260807 476176
rect 259564 476172 259570 476174
rect 260741 476171 260807 476174
rect 261702 476172 261708 476236
rect 261772 476234 261778 476236
rect 262857 476234 262923 476237
rect 261772 476232 262923 476234
rect 261772 476176 262862 476232
rect 262918 476176 262923 476232
rect 261772 476174 262923 476176
rect 261772 476172 261778 476174
rect 262857 476171 262923 476174
rect 265382 476172 265388 476236
rect 265452 476234 265458 476236
rect 266261 476234 266327 476237
rect 265452 476232 266327 476234
rect 265452 476176 266266 476232
rect 266322 476176 266327 476232
rect 265452 476174 266327 476176
rect 265452 476172 265458 476174
rect 266261 476171 266327 476174
rect 266486 476172 266492 476236
rect 266556 476234 266562 476236
rect 267641 476234 267707 476237
rect 266556 476232 267707 476234
rect 266556 476176 267646 476232
rect 267702 476176 267707 476232
rect 266556 476174 267707 476176
rect 266556 476172 266562 476174
rect 267641 476171 267707 476174
rect 268694 476172 268700 476236
rect 268764 476234 268770 476236
rect 269021 476234 269087 476237
rect 268764 476232 269087 476234
rect 268764 476176 269026 476232
rect 269082 476176 269087 476232
rect 268764 476174 269087 476176
rect 268764 476172 268770 476174
rect 269021 476171 269087 476174
rect 269798 476172 269804 476236
rect 269868 476234 269874 476236
rect 270401 476234 270467 476237
rect 269868 476232 270467 476234
rect 269868 476176 270406 476232
rect 270462 476176 270467 476232
rect 269868 476174 270467 476176
rect 269868 476172 269874 476174
rect 270401 476171 270467 476174
rect 271270 476172 271276 476236
rect 271340 476234 271346 476236
rect 271781 476234 271847 476237
rect 271340 476232 271847 476234
rect 271340 476176 271786 476232
rect 271842 476176 271847 476232
rect 271340 476174 271847 476176
rect 271340 476172 271346 476174
rect 271781 476171 271847 476174
rect 272190 476172 272196 476236
rect 272260 476234 272266 476236
rect 273161 476234 273227 476237
rect 272260 476232 273227 476234
rect 272260 476176 273166 476232
rect 273222 476176 273227 476232
rect 272260 476174 273227 476176
rect 272260 476172 272266 476174
rect 273161 476171 273227 476174
rect 273294 476172 273300 476236
rect 273364 476234 273370 476236
rect 274541 476234 274607 476237
rect 275921 476236 275987 476237
rect 273364 476232 274607 476234
rect 273364 476176 274546 476232
rect 274602 476176 274607 476232
rect 273364 476174 274607 476176
rect 273364 476172 273370 476174
rect 274541 476171 274607 476174
rect 275870 476172 275876 476236
rect 275940 476234 275987 476236
rect 275940 476232 276032 476234
rect 275982 476176 276032 476232
rect 275940 476174 276032 476176
rect 275940 476172 275987 476174
rect 276974 476172 276980 476236
rect 277044 476234 277050 476236
rect 277301 476234 277367 476237
rect 277044 476232 277367 476234
rect 277044 476176 277306 476232
rect 277362 476176 277367 476232
rect 277044 476174 277367 476176
rect 277044 476172 277050 476174
rect 275921 476171 275987 476172
rect 277301 476171 277367 476174
rect 278078 476172 278084 476236
rect 278148 476234 278154 476236
rect 278681 476234 278747 476237
rect 278148 476232 278747 476234
rect 278148 476176 278686 476232
rect 278742 476176 278747 476232
rect 278148 476174 278747 476176
rect 278148 476172 278154 476174
rect 278681 476171 278747 476174
rect 279182 476172 279188 476236
rect 279252 476234 279258 476236
rect 280061 476234 280127 476237
rect 279252 476232 280127 476234
rect 279252 476176 280066 476232
rect 280122 476176 280127 476232
rect 279252 476174 280127 476176
rect 279252 476172 279258 476174
rect 280061 476171 280127 476174
rect 280245 476234 280311 476237
rect 280838 476234 280844 476236
rect 280245 476232 280844 476234
rect 280245 476176 280250 476232
rect 280306 476176 280844 476232
rect 280245 476174 280844 476176
rect 280245 476171 280311 476174
rect 280838 476172 280844 476174
rect 280908 476172 280914 476236
rect 283005 476234 283071 476237
rect 283414 476234 283420 476236
rect 283005 476232 283420 476234
rect 283005 476176 283010 476232
rect 283066 476176 283420 476232
rect 283005 476174 283420 476176
rect 283005 476171 283071 476174
rect 283414 476172 283420 476174
rect 283484 476172 283490 476236
rect 285765 476234 285831 476237
rect 285990 476234 285996 476236
rect 285765 476232 285996 476234
rect 285765 476176 285770 476232
rect 285826 476176 285996 476232
rect 285765 476174 285996 476176
rect 285765 476171 285831 476174
rect 285990 476172 285996 476174
rect 286060 476172 286066 476236
rect 287053 476234 287119 476237
rect 288198 476234 288204 476236
rect 287053 476232 288204 476234
rect 287053 476176 287058 476232
rect 287114 476176 288204 476232
rect 287053 476174 288204 476176
rect 287053 476171 287119 476174
rect 288198 476172 288204 476174
rect 288268 476172 288274 476236
rect 289905 476234 289971 476237
rect 290958 476234 290964 476236
rect 289905 476232 290964 476234
rect 289905 476176 289910 476232
rect 289966 476176 290964 476232
rect 289905 476174 290964 476176
rect 289905 476171 289971 476174
rect 290958 476172 290964 476174
rect 291028 476172 291034 476236
rect 292573 476234 292639 476237
rect 293350 476234 293356 476236
rect 292573 476232 293356 476234
rect 292573 476176 292578 476232
rect 292634 476176 293356 476232
rect 292573 476174 293356 476176
rect 292573 476171 292639 476174
rect 293350 476172 293356 476174
rect 293420 476172 293426 476236
rect 295425 476234 295491 476237
rect 295926 476234 295932 476236
rect 295425 476232 295932 476234
rect 295425 476176 295430 476232
rect 295486 476176 295932 476232
rect 295425 476174 295932 476176
rect 295425 476171 295491 476174
rect 295926 476172 295932 476174
rect 295996 476172 296002 476236
rect 298185 476234 298251 476237
rect 300945 476236 301011 476237
rect 298502 476234 298508 476236
rect 298185 476232 298508 476234
rect 298185 476176 298190 476232
rect 298246 476176 298508 476232
rect 298185 476174 298508 476176
rect 298185 476171 298251 476174
rect 298502 476172 298508 476174
rect 298572 476172 298578 476236
rect 300894 476172 300900 476236
rect 300964 476234 301011 476236
rect 300964 476232 301056 476234
rect 301006 476176 301056 476232
rect 300964 476174 301056 476176
rect 300964 476172 301011 476174
rect 300945 476171 301011 476172
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 583520 471324 584960 471564
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 2865 449578 2931 449581
rect -960 449576 2931 449578
rect -960 449520 2870 449576
rect 2926 449520 2931 449576
rect -960 449518 2931 449520
rect -960 449428 480 449518
rect 2865 449515 2931 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580349 431626 580415 431629
rect 583520 431626 584960 431716
rect 580349 431624 584960 431626
rect 580349 431568 580354 431624
rect 580410 431568 584960 431624
rect 580349 431566 584960 431568
rect 580349 431563 580415 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 583520 404820 584960 405060
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3049 371378 3115 371381
rect -960 371376 3115 371378
rect -960 371320 3054 371376
rect 3110 371320 3115 371376
rect -960 371318 3115 371320
rect -960 371228 480 371318
rect 3049 371315 3115 371318
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 583520 311932 584960 312172
rect 282678 309028 282684 309092
rect 282748 309090 282754 309092
rect 298093 309090 298159 309093
rect 282748 309088 298159 309090
rect 282748 309032 298098 309088
rect 298154 309032 298159 309088
rect 282748 309030 298159 309032
rect 282748 309028 282754 309030
rect 298093 309027 298159 309030
rect 283414 308892 283420 308956
rect 283484 308954 283490 308956
rect 348325 308954 348391 308957
rect 283484 308952 348391 308954
rect 283484 308896 348330 308952
rect 348386 308896 348391 308952
rect 283484 308894 348391 308896
rect 283484 308892 283490 308894
rect 348325 308891 348391 308894
rect 282126 308756 282132 308820
rect 282196 308818 282202 308820
rect 349613 308818 349679 308821
rect 282196 308816 349679 308818
rect 282196 308760 349618 308816
rect 349674 308760 349679 308816
rect 282196 308758 349679 308760
rect 282196 308756 282202 308758
rect 349613 308755 349679 308758
rect 250989 308682 251055 308685
rect 347037 308682 347103 308685
rect 250989 308680 347103 308682
rect 250989 308624 250994 308680
rect 251050 308624 347042 308680
rect 347098 308624 347103 308680
rect 250989 308622 347103 308624
rect 250989 308619 251055 308622
rect 347037 308619 347103 308622
rect 284702 308484 284708 308548
rect 284772 308546 284778 308548
rect 352281 308546 352347 308549
rect 284772 308544 352347 308546
rect 284772 308488 352286 308544
rect 352342 308488 352347 308544
rect 284772 308486 352347 308488
rect 284772 308484 284778 308486
rect 352281 308483 352347 308486
rect 238201 308410 238267 308413
rect 337929 308410 337995 308413
rect 238201 308408 337995 308410
rect 238201 308352 238206 308408
rect 238262 308352 337934 308408
rect 337990 308352 337995 308408
rect 238201 308350 337995 308352
rect 238201 308347 238267 308350
rect 337929 308347 337995 308350
rect 296989 308274 297055 308277
rect 297950 308274 297956 308276
rect 296989 308272 297956 308274
rect 296989 308216 296994 308272
rect 297050 308216 297956 308272
rect 296989 308214 297956 308216
rect 296989 308211 297055 308214
rect 297950 308212 297956 308214
rect 298020 308212 298026 308276
rect 297398 308076 297404 308140
rect 297468 308138 297474 308140
rect 297909 308138 297975 308141
rect 297468 308136 297975 308138
rect 297468 308080 297914 308136
rect 297970 308080 297975 308136
rect 297468 308078 297975 308080
rect 297468 308076 297474 308078
rect 297909 308075 297975 308078
rect 277342 307940 277348 308004
rect 277412 308002 277418 308004
rect 277485 308002 277551 308005
rect 277412 308000 277551 308002
rect 277412 307944 277490 308000
rect 277546 307944 277551 308000
rect 277412 307942 277551 307944
rect 277412 307940 277418 307942
rect 277485 307939 277551 307942
rect 297265 308002 297331 308005
rect 297582 308002 297588 308004
rect 297265 308000 297588 308002
rect 297265 307944 297270 308000
rect 297326 307944 297588 308000
rect 297265 307942 297588 307944
rect 297265 307939 297331 307942
rect 297582 307940 297588 307942
rect 297652 307940 297658 308004
rect 298318 307940 298324 308004
rect 298388 308002 298394 308004
rect 299197 308002 299263 308005
rect 298388 308000 299263 308002
rect 298388 307944 299202 308000
rect 299258 307944 299263 308000
rect 298388 307942 299263 307944
rect 298388 307940 298394 307942
rect 299197 307939 299263 307942
rect 277526 307804 277532 307868
rect 277596 307866 277602 307868
rect 277669 307866 277735 307869
rect 277596 307864 277735 307866
rect 277596 307808 277674 307864
rect 277730 307808 277735 307864
rect 277596 307806 277735 307808
rect 277596 307804 277602 307806
rect 277669 307803 277735 307806
rect 278773 307868 278839 307869
rect 278773 307864 278820 307868
rect 278884 307866 278890 307868
rect 278773 307808 278778 307864
rect 278773 307804 278820 307808
rect 278884 307806 278930 307866
rect 278884 307804 278890 307806
rect 278998 307804 279004 307868
rect 279068 307866 279074 307868
rect 279233 307866 279299 307869
rect 279068 307864 279299 307866
rect 279068 307808 279238 307864
rect 279294 307808 279299 307864
rect 279068 307806 279299 307808
rect 279068 307804 279074 307806
rect 278773 307803 278839 307804
rect 279233 307803 279299 307806
rect 284886 307804 284892 307868
rect 284956 307866 284962 307868
rect 285489 307866 285555 307869
rect 284956 307864 285555 307866
rect 284956 307808 285494 307864
rect 285550 307808 285555 307864
rect 284956 307806 285555 307808
rect 284956 307804 284962 307806
rect 285489 307803 285555 307806
rect 296478 307804 296484 307868
rect 296548 307866 296554 307868
rect 296621 307866 296687 307869
rect 296548 307864 296687 307866
rect 296548 307808 296626 307864
rect 296682 307808 296687 307864
rect 296548 307806 296687 307808
rect 296548 307804 296554 307806
rect 296621 307803 296687 307806
rect 297633 307866 297699 307869
rect 297766 307866 297772 307868
rect 297633 307864 297772 307866
rect 297633 307808 297638 307864
rect 297694 307808 297772 307864
rect 297633 307806 297772 307808
rect 297633 307803 297699 307806
rect 297766 307804 297772 307806
rect 297836 307804 297842 307868
rect 298502 307804 298508 307868
rect 298572 307866 298578 307868
rect 299013 307866 299079 307869
rect 298572 307864 299079 307866
rect 298572 307808 299018 307864
rect 299074 307808 299079 307864
rect 298572 307806 299079 307808
rect 298572 307804 298578 307806
rect 299013 307803 299079 307806
rect 316125 307866 316191 307869
rect 318149 307866 318215 307869
rect 316125 307864 318215 307866
rect 316125 307808 316130 307864
rect 316186 307808 318154 307864
rect 318210 307808 318215 307864
rect 316125 307806 318215 307808
rect 316125 307803 316191 307806
rect 318149 307803 318215 307806
rect 241973 306370 242039 306373
rect 318977 306370 319043 306373
rect 320081 306370 320147 306373
rect 241973 306368 242082 306370
rect -960 306234 480 306324
rect 241973 306312 241978 306368
rect 242034 306312 242082 306368
rect 241973 306307 242082 306312
rect 318977 306368 320147 306370
rect 318977 306312 318982 306368
rect 319038 306312 320086 306368
rect 320142 306312 320147 306368
rect 318977 306310 320147 306312
rect 318977 306307 319043 306310
rect 320081 306307 320147 306310
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 242022 306101 242082 306307
rect 279325 306234 279391 306237
rect 280061 306234 280127 306237
rect 279325 306232 280127 306234
rect 279325 306176 279330 306232
rect 279386 306176 280066 306232
rect 280122 306176 280127 306232
rect 279325 306174 280127 306176
rect 279325 306171 279391 306174
rect 280061 306171 280127 306174
rect 283782 306172 283788 306236
rect 283852 306234 283858 306236
rect 338941 306234 339007 306237
rect 283852 306232 339007 306234
rect 283852 306176 338946 306232
rect 339002 306176 339007 306232
rect 283852 306174 339007 306176
rect 283852 306172 283858 306174
rect 338941 306171 339007 306174
rect 241973 306096 242082 306101
rect 241973 306040 241978 306096
rect 242034 306040 242082 306096
rect 241973 306038 242082 306040
rect 270493 306098 270559 306101
rect 270861 306098 270927 306101
rect 270493 306096 270927 306098
rect 270493 306040 270498 306096
rect 270554 306040 270866 306096
rect 270922 306040 270927 306096
rect 270493 306038 270927 306040
rect 241973 306035 242039 306038
rect 270493 306035 270559 306038
rect 270861 306035 270927 306038
rect 283598 306036 283604 306100
rect 283668 306098 283674 306100
rect 353385 306098 353451 306101
rect 283668 306096 353451 306098
rect 283668 306040 353390 306096
rect 353446 306040 353451 306096
rect 283668 306038 353451 306040
rect 283668 306036 283674 306038
rect 353385 306035 353451 306038
rect 312629 305962 312695 305965
rect 442257 305962 442323 305965
rect 312629 305960 442323 305962
rect 312629 305904 312634 305960
rect 312690 305904 442262 305960
rect 442318 305904 442323 305960
rect 312629 305902 442323 305904
rect 312629 305899 312695 305902
rect 442257 305899 442323 305902
rect 320081 305826 320147 305829
rect 476757 305826 476823 305829
rect 320081 305824 476823 305826
rect 320081 305768 320086 305824
rect 320142 305768 476762 305824
rect 476818 305768 476823 305824
rect 320081 305766 476823 305768
rect 320081 305763 320147 305766
rect 476757 305763 476823 305766
rect 324221 305690 324287 305693
rect 511993 305690 512059 305693
rect 324221 305688 512059 305690
rect 324221 305632 324226 305688
rect 324282 305632 511998 305688
rect 512054 305632 512059 305688
rect 324221 305630 512059 305632
rect 324221 305627 324287 305630
rect 511993 305627 512059 305630
rect 324405 305554 324471 305557
rect 324589 305554 324655 305557
rect 324405 305552 324655 305554
rect 324405 305496 324410 305552
rect 324466 305496 324594 305552
rect 324650 305496 324655 305552
rect 324405 305494 324655 305496
rect 324405 305491 324471 305494
rect 324589 305491 324655 305494
rect 331397 305554 331463 305557
rect 331673 305554 331739 305557
rect 331397 305552 331739 305554
rect 331397 305496 331402 305552
rect 331458 305496 331678 305552
rect 331734 305496 331739 305552
rect 331397 305494 331739 305496
rect 331397 305491 331463 305494
rect 331673 305491 331739 305494
rect 275318 303316 275324 303380
rect 275388 303378 275394 303380
rect 340045 303378 340111 303381
rect 275388 303376 340111 303378
rect 275388 303320 340050 303376
rect 340106 303320 340111 303376
rect 275388 303318 340111 303320
rect 275388 303316 275394 303318
rect 340045 303315 340111 303318
rect 275134 303180 275140 303244
rect 275204 303242 275210 303244
rect 341057 303242 341123 303245
rect 275204 303240 341123 303242
rect 275204 303184 341062 303240
rect 341118 303184 341123 303240
rect 275204 303182 341123 303184
rect 275204 303180 275210 303182
rect 341057 303179 341123 303182
rect 272609 303106 272675 303109
rect 342437 303106 342503 303109
rect 272609 303104 342503 303106
rect 272609 303048 272614 303104
rect 272670 303048 342442 303104
rect 342498 303048 342503 303104
rect 272609 303046 342503 303048
rect 272609 303043 272675 303046
rect 342437 303043 342503 303046
rect 311617 302970 311683 302973
rect 439446 302970 439452 302972
rect 311617 302968 439452 302970
rect 311617 302912 311622 302968
rect 311678 302912 439452 302968
rect 311617 302910 439452 302912
rect 311617 302907 311683 302910
rect 439446 302908 439452 302910
rect 439516 302908 439522 302972
rect 321093 302834 321159 302837
rect 489913 302834 489979 302837
rect 321093 302832 489979 302834
rect 321093 302776 321098 302832
rect 321154 302776 489918 302832
rect 489974 302776 489979 302832
rect 321093 302774 489979 302776
rect 321093 302771 321159 302774
rect 489913 302771 489979 302774
rect 279693 300658 279759 300661
rect 352649 300658 352715 300661
rect 279693 300656 352715 300658
rect 279693 300600 279698 300656
rect 279754 300600 352654 300656
rect 352710 300600 352715 300656
rect 279693 300598 352715 300600
rect 279693 300595 279759 300598
rect 352649 300595 352715 300598
rect 281349 300522 281415 300525
rect 356421 300522 356487 300525
rect 281349 300520 356487 300522
rect 281349 300464 281354 300520
rect 281410 300464 356426 300520
rect 356482 300464 356487 300520
rect 281349 300462 356487 300464
rect 281349 300459 281415 300462
rect 356421 300459 356487 300462
rect 279785 300386 279851 300389
rect 355777 300386 355843 300389
rect 279785 300384 355843 300386
rect 279785 300328 279790 300384
rect 279846 300328 355782 300384
rect 355838 300328 355843 300384
rect 279785 300326 355843 300328
rect 279785 300323 279851 300326
rect 355777 300323 355843 300326
rect 278681 300250 278747 300253
rect 359181 300250 359247 300253
rect 278681 300248 359247 300250
rect 278681 300192 278686 300248
rect 278742 300192 359186 300248
rect 359242 300192 359247 300248
rect 278681 300190 359247 300192
rect 278681 300187 278747 300190
rect 359181 300187 359247 300190
rect 321921 300114 321987 300117
rect 498285 300114 498351 300117
rect 321921 300112 498351 300114
rect 321921 300056 321926 300112
rect 321982 300056 498290 300112
rect 498346 300056 498351 300112
rect 321921 300054 498351 300056
rect 321921 300051 321987 300054
rect 498285 300051 498351 300054
rect 310973 298754 311039 298757
rect 439078 298754 439084 298756
rect 310973 298752 439084 298754
rect 310973 298696 310978 298752
rect 311034 298696 439084 298752
rect 310973 298694 439084 298696
rect 310973 298691 311039 298694
rect 439078 298692 439084 298694
rect 439148 298692 439154 298756
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 310881 287738 310947 287741
rect 437422 287738 437428 287740
rect 310881 287736 437428 287738
rect 310881 287680 310886 287736
rect 310942 287680 437428 287736
rect 310881 287678 437428 287680
rect 310881 287675 310947 287678
rect 437422 287676 437428 287678
rect 437492 287676 437498 287740
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 287646 248100 287652 248164
rect 287716 248162 287722 248164
rect 299841 248162 299907 248165
rect 287716 248160 299907 248162
rect 287716 248104 299846 248160
rect 299902 248104 299907 248160
rect 287716 248102 299907 248104
rect 287716 248100 287722 248102
rect 299841 248099 299907 248102
rect 286910 247964 286916 248028
rect 286980 248026 286986 248028
rect 299933 248026 299999 248029
rect 286980 248024 299999 248026
rect 286980 247968 299938 248024
rect 299994 247968 299999 248024
rect 286980 247966 299999 247968
rect 286980 247964 286986 247966
rect 299933 247963 299999 247966
rect 300669 248026 300735 248029
rect 305269 248026 305335 248029
rect 300669 248024 305335 248026
rect 300669 247968 300674 248024
rect 300730 247968 305274 248024
rect 305330 247968 305335 248024
rect 300669 247966 305335 247968
rect 300669 247963 300735 247966
rect 305269 247963 305335 247966
rect 289486 247828 289492 247892
rect 289556 247890 289562 247892
rect 302785 247890 302851 247893
rect 289556 247888 302851 247890
rect 289556 247832 302790 247888
rect 302846 247832 302851 247888
rect 289556 247830 302851 247832
rect 289556 247828 289562 247830
rect 302785 247827 302851 247830
rect 288198 247692 288204 247756
rect 288268 247754 288274 247756
rect 302601 247754 302667 247757
rect 288268 247752 302667 247754
rect 288268 247696 302606 247752
rect 302662 247696 302667 247752
rect 288268 247694 302667 247696
rect 288268 247692 288274 247694
rect 302601 247691 302667 247694
rect 286542 247556 286548 247620
rect 286612 247618 286618 247620
rect 301221 247618 301287 247621
rect 286612 247616 301287 247618
rect 286612 247560 301226 247616
rect 301282 247560 301287 247616
rect 286612 247558 301287 247560
rect 286612 247556 286618 247558
rect 301221 247555 301287 247558
rect 308121 247618 308187 247621
rect 437606 247618 437612 247620
rect 308121 247616 437612 247618
rect 308121 247560 308126 247616
rect 308182 247560 437612 247616
rect 308121 247558 437612 247560
rect 308121 247555 308187 247558
rect 437606 247556 437612 247558
rect 437676 247556 437682 247620
rect 295190 247420 295196 247484
rect 295260 247482 295266 247484
rect 302693 247482 302759 247485
rect 295260 247480 302759 247482
rect 295260 247424 302698 247480
rect 302754 247424 302759 247480
rect 295260 247422 302759 247424
rect 295260 247420 295266 247422
rect 302693 247419 302759 247422
rect 293534 247284 293540 247348
rect 293604 247346 293610 247348
rect 301313 247346 301379 247349
rect 293604 247344 301379 247346
rect 293604 247288 301318 247344
rect 301374 247288 301379 247344
rect 293604 247286 301379 247288
rect 293604 247284 293610 247286
rect 301313 247283 301379 247286
rect 286777 247076 286843 247077
rect 287881 247076 287947 247077
rect 288065 247076 288131 247077
rect 288985 247076 289051 247077
rect 289169 247076 289235 247077
rect 290641 247076 290707 247077
rect 286726 247074 286732 247076
rect 286686 247014 286732 247074
rect 286796 247072 286843 247076
rect 287830 247074 287836 247076
rect 286838 247016 286843 247072
rect 286726 247012 286732 247014
rect 286796 247012 286843 247016
rect 287790 247014 287836 247074
rect 287900 247072 287947 247076
rect 287942 247016 287947 247072
rect 287830 247012 287836 247014
rect 287900 247012 287947 247016
rect 288014 247012 288020 247076
rect 288084 247074 288131 247076
rect 288934 247074 288940 247076
rect 288084 247072 288176 247074
rect 288126 247016 288176 247072
rect 288084 247014 288176 247016
rect 288894 247014 288940 247074
rect 289004 247072 289051 247076
rect 289046 247016 289051 247072
rect 288084 247012 288131 247014
rect 288934 247012 288940 247014
rect 289004 247012 289051 247016
rect 289118 247012 289124 247076
rect 289188 247074 289235 247076
rect 290590 247074 290596 247076
rect 289188 247072 289280 247074
rect 289230 247016 289280 247072
rect 289188 247014 289280 247016
rect 290550 247014 290596 247074
rect 290660 247072 290707 247076
rect 290702 247016 290707 247072
rect 289188 247012 289235 247014
rect 290590 247012 290596 247014
rect 290660 247012 290707 247016
rect 292246 247012 292252 247076
rect 292316 247074 292322 247076
rect 292389 247074 292455 247077
rect 292316 247072 292455 247074
rect 292316 247016 292394 247072
rect 292450 247016 292455 247072
rect 292316 247014 292455 247016
rect 292316 247012 292322 247014
rect 286777 247011 286843 247012
rect 287881 247011 287947 247012
rect 288065 247011 288131 247012
rect 288985 247011 289051 247012
rect 289169 247011 289235 247012
rect 290641 247011 290707 247012
rect 292389 247011 292455 247014
rect 285070 246196 285076 246260
rect 285140 246258 285146 246260
rect 296805 246258 296871 246261
rect 285140 246256 296871 246258
rect 285140 246200 296810 246256
rect 296866 246200 296871 246256
rect 285140 246198 296871 246200
rect 285140 246196 285146 246198
rect 296805 246195 296871 246198
rect 299289 245578 299355 245581
rect 306557 245578 306623 245581
rect 299289 245576 306623 245578
rect 299289 245520 299294 245576
rect 299350 245520 306562 245576
rect 306618 245520 306623 245576
rect 299289 245518 306623 245520
rect 299289 245515 299355 245518
rect 306557 245515 306623 245518
rect 295926 245380 295932 245444
rect 295996 245442 296002 245444
rect 302325 245442 302391 245445
rect 295996 245440 302391 245442
rect 295996 245384 302330 245440
rect 302386 245384 302391 245440
rect 583520 245428 584960 245668
rect 295996 245382 302391 245384
rect 295996 245380 296002 245382
rect 302325 245379 302391 245382
rect 292430 245244 292436 245308
rect 292500 245306 292506 245308
rect 300945 245306 301011 245309
rect 292500 245304 301011 245306
rect 292500 245248 300950 245304
rect 301006 245248 301011 245304
rect 292500 245246 301011 245248
rect 292500 245244 292506 245246
rect 300945 245243 301011 245246
rect 309225 245306 309291 245309
rect 437790 245306 437796 245308
rect 309225 245304 437796 245306
rect 309225 245248 309230 245304
rect 309286 245248 437796 245304
rect 309225 245246 437796 245248
rect 309225 245243 309291 245246
rect 437790 245244 437796 245246
rect 437860 245244 437866 245308
rect 290774 245108 290780 245172
rect 290844 245170 290850 245172
rect 291009 245170 291075 245173
rect 290844 245168 291075 245170
rect 290844 245112 291014 245168
rect 291070 245112 291075 245168
rect 290844 245110 291075 245112
rect 290844 245108 290850 245110
rect 291009 245107 291075 245110
rect 293718 245108 293724 245172
rect 293788 245170 293794 245172
rect 302417 245170 302483 245173
rect 293788 245168 302483 245170
rect 293788 245112 302422 245168
rect 302478 245112 302483 245168
rect 293788 245110 302483 245112
rect 293788 245108 293794 245110
rect 302417 245107 302483 245110
rect 324313 245170 324379 245173
rect 516133 245170 516199 245173
rect 324313 245168 516199 245170
rect 324313 245112 324318 245168
rect 324374 245112 516138 245168
rect 516194 245112 516199 245168
rect 324313 245110 516199 245112
rect 324313 245107 324379 245110
rect 516133 245107 516199 245110
rect 289302 244972 289308 245036
rect 289372 245034 289378 245036
rect 302509 245034 302575 245037
rect 289372 245032 302575 245034
rect 289372 244976 302514 245032
rect 302570 244976 302575 245032
rect 289372 244974 302575 244976
rect 289372 244972 289378 244974
rect 302509 244971 302575 244974
rect 325693 245034 325759 245037
rect 523125 245034 523191 245037
rect 325693 245032 523191 245034
rect 325693 244976 325698 245032
rect 325754 244976 523130 245032
rect 523186 244976 523191 245032
rect 325693 244974 523191 244976
rect 325693 244971 325759 244974
rect 523125 244971 523191 244974
rect 282494 244836 282500 244900
rect 282564 244898 282570 244900
rect 296713 244898 296779 244901
rect 282564 244896 296779 244898
rect 282564 244840 296718 244896
rect 296774 244840 296779 244896
rect 282564 244838 296779 244840
rect 282564 244836 282570 244838
rect 296713 244835 296779 244838
rect 327073 244898 327139 244901
rect 531405 244898 531471 244901
rect 327073 244896 531471 244898
rect 327073 244840 327078 244896
rect 327134 244840 531410 244896
rect 531466 244840 531471 244896
rect 327073 244838 531471 244840
rect 327073 244835 327139 244838
rect 531405 244835 531471 244838
rect 295006 244700 295012 244764
rect 295076 244762 295082 244764
rect 295241 244762 295307 244765
rect 295076 244760 295307 244762
rect 295076 244704 295246 244760
rect 295302 244704 295307 244760
rect 295076 244702 295307 244704
rect 295076 244700 295082 244702
rect 295241 244699 295307 244702
rect 296110 244700 296116 244764
rect 296180 244762 296186 244764
rect 301037 244762 301103 244765
rect 296180 244760 301103 244762
rect 296180 244704 301042 244760
rect 301098 244704 301103 244760
rect 296180 244702 301103 244704
rect 296180 244700 296186 244702
rect 301037 244699 301103 244702
rect 296294 244564 296300 244628
rect 296364 244626 296370 244628
rect 299749 244626 299815 244629
rect 296364 244624 299815 244626
rect 296364 244568 299754 244624
rect 299810 244568 299815 244624
rect 296364 244566 299815 244568
rect 296364 244564 296370 244566
rect 299749 244563 299815 244566
rect 293166 244428 293172 244492
rect 293236 244490 293242 244492
rect 293401 244490 293467 244493
rect 293236 244488 293467 244490
rect 293236 244432 293406 244488
rect 293462 244432 293467 244488
rect 293236 244430 293467 244432
rect 293236 244428 293242 244430
rect 293401 244427 293467 244430
rect 291745 244356 291811 244357
rect 291694 244354 291700 244356
rect 291654 244294 291700 244354
rect 291764 244352 291811 244356
rect 291806 244296 291811 244352
rect 291694 244292 291700 244294
rect 291764 244292 291811 244296
rect 291878 244292 291884 244356
rect 291948 244354 291954 244356
rect 292205 244354 292271 244357
rect 291948 244352 292271 244354
rect 291948 244296 292210 244352
rect 292266 244296 292271 244352
rect 291948 244294 292271 244296
rect 291948 244292 291954 244294
rect 291745 244291 291811 244292
rect 292205 244291 292271 244294
rect 293350 244292 293356 244356
rect 293420 244354 293426 244356
rect 293677 244354 293743 244357
rect 293420 244352 293743 244354
rect 293420 244296 293682 244352
rect 293738 244296 293743 244352
rect 293420 244294 293743 244296
rect 293420 244292 293426 244294
rect 293677 244291 293743 244294
rect 298134 244292 298140 244356
rect 298204 244354 298210 244356
rect 298369 244354 298435 244357
rect 298737 244356 298803 244357
rect 298686 244354 298692 244356
rect 298204 244352 298435 244354
rect 298204 244296 298374 244352
rect 298430 244296 298435 244352
rect 298204 244294 298435 244296
rect 298646 244294 298692 244354
rect 298756 244352 298803 244356
rect 298798 244296 298803 244352
rect 298204 244292 298210 244294
rect 298369 244291 298435 244294
rect 298686 244292 298692 244294
rect 298756 244292 298803 244296
rect 298737 244291 298803 244292
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 97717 196890 97783 196893
rect 99422 196890 100004 196924
rect 97717 196888 100004 196890
rect 97717 196832 97722 196888
rect 97778 196864 100004 196888
rect 298921 196890 298987 196893
rect 299430 196890 300012 196924
rect 298921 196888 300012 196890
rect 97778 196832 99482 196864
rect 97717 196830 99482 196832
rect 298921 196832 298926 196888
rect 298982 196864 300012 196888
rect 298982 196832 299490 196864
rect 298921 196830 299490 196832
rect 97717 196827 97783 196830
rect 298921 196827 298987 196830
rect 291878 196012 291884 196076
rect 291948 196074 291954 196076
rect 292113 196074 292179 196077
rect 291948 196072 292179 196074
rect 291948 196016 292118 196072
rect 292174 196016 292179 196072
rect 291948 196014 292179 196016
rect 291948 196012 291954 196014
rect 292113 196011 292179 196014
rect 97809 195938 97875 195941
rect 99422 195938 100004 195972
rect 97809 195936 100004 195938
rect 97809 195880 97814 195936
rect 97870 195912 100004 195936
rect 297265 195938 297331 195941
rect 299430 195938 300012 195972
rect 297265 195936 300012 195938
rect 97870 195880 99482 195912
rect 97809 195878 99482 195880
rect 297265 195880 297270 195936
rect 297326 195912 300012 195936
rect 297326 195880 299490 195912
rect 297265 195878 299490 195880
rect 97809 195875 97875 195878
rect 297265 195875 297331 195878
rect 97809 193762 97875 193765
rect 99422 193762 100004 193796
rect 97809 193760 100004 193762
rect 97809 193704 97814 193760
rect 97870 193736 100004 193760
rect 299105 193762 299171 193765
rect 299430 193762 300012 193796
rect 299105 193760 300012 193762
rect 97870 193704 99482 193736
rect 97809 193702 99482 193704
rect 299105 193704 299110 193760
rect 299166 193736 300012 193760
rect 299166 193704 299490 193736
rect 299105 193702 299490 193704
rect 97809 193699 97875 193702
rect 299105 193699 299171 193702
rect 97533 192810 97599 192813
rect 99422 192810 100004 192844
rect 97533 192808 100004 192810
rect 97533 192752 97538 192808
rect 97594 192784 100004 192808
rect 297357 192810 297423 192813
rect 299430 192810 300012 192844
rect 297357 192808 300012 192810
rect 97594 192752 99482 192784
rect 97533 192750 99482 192752
rect 297357 192752 297362 192808
rect 297418 192784 300012 192808
rect 297418 192752 299490 192784
rect 297357 192750 299490 192752
rect 97533 192747 97599 192750
rect 297357 192747 297423 192750
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect 297265 191722 297331 191725
rect 297449 191722 297515 191725
rect 297265 191720 297515 191722
rect 297265 191664 297270 191720
rect 297326 191664 297454 191720
rect 297510 191664 297515 191720
rect 297265 191662 297515 191664
rect 297265 191659 297331 191662
rect 297449 191659 297515 191662
rect 97625 191042 97691 191045
rect 99422 191042 100004 191076
rect 97625 191040 100004 191042
rect 97625 190984 97630 191040
rect 97686 191016 100004 191040
rect 297265 191042 297331 191045
rect 299430 191042 300012 191076
rect 297265 191040 300012 191042
rect 97686 190984 99482 191016
rect 97625 190982 99482 190984
rect 297265 190984 297270 191040
rect 297326 191016 300012 191040
rect 297326 190984 299490 191016
rect 297265 190982 299490 190984
rect 97625 190979 97691 190982
rect 297265 190979 297331 190982
rect 97717 189954 97783 189957
rect 99422 189954 100004 189988
rect 97717 189952 100004 189954
rect 97717 189896 97722 189952
rect 97778 189928 100004 189952
rect 297081 189954 297147 189957
rect 299430 189954 300012 189988
rect 297081 189952 300012 189954
rect 97778 189896 99482 189928
rect 97717 189894 99482 189896
rect 297081 189896 297086 189952
rect 297142 189928 300012 189952
rect 297142 189896 299490 189928
rect 297081 189894 299490 189896
rect 97717 189891 97783 189894
rect 297081 189891 297147 189894
rect 297081 189138 297147 189141
rect 297449 189138 297515 189141
rect 297081 189136 297515 189138
rect 297081 189080 297086 189136
rect 297142 189080 297454 189136
rect 297510 189080 297515 189136
rect 297081 189078 297515 189080
rect 297081 189075 297147 189078
rect 297449 189075 297515 189078
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 97901 188186 97967 188189
rect 99422 188186 100004 188220
rect 97901 188184 100004 188186
rect 97901 188128 97906 188184
rect 97962 188160 100004 188184
rect 298737 188186 298803 188189
rect 299430 188186 300012 188220
rect 298737 188184 300012 188186
rect 97962 188128 99482 188160
rect 97901 188126 99482 188128
rect 298737 188128 298742 188184
rect 298798 188160 300012 188184
rect 298798 188128 299490 188160
rect 298737 188126 299490 188128
rect 97901 188123 97967 188126
rect 298737 188123 298803 188126
rect 298134 187716 298140 187780
rect 298204 187778 298210 187780
rect 299105 187778 299171 187781
rect 298204 187776 299171 187778
rect 298204 187720 299110 187776
rect 299166 187720 299171 187776
rect 298204 187718 299171 187720
rect 298204 187716 298210 187718
rect 299105 187715 299171 187718
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 97901 169962 97967 169965
rect 99422 169962 100004 169996
rect 97901 169960 100004 169962
rect 97901 169904 97906 169960
rect 97962 169936 100004 169960
rect 297173 169962 297239 169965
rect 299430 169962 300012 169996
rect 297173 169960 300012 169962
rect 97962 169904 99482 169936
rect 97901 169902 99482 169904
rect 297173 169904 297178 169960
rect 297234 169936 300012 169960
rect 297234 169904 299490 169936
rect 297173 169902 299490 169904
rect 97901 169899 97967 169902
rect 297173 169899 297239 169902
rect 97441 168330 97507 168333
rect 99422 168330 100004 168364
rect 97441 168328 100004 168330
rect 97441 168272 97446 168328
rect 97502 168304 100004 168328
rect 297725 168330 297791 168333
rect 299430 168330 300012 168364
rect 297725 168328 300012 168330
rect 97502 168272 99482 168304
rect 97441 168270 99482 168272
rect 297725 168272 297730 168328
rect 297786 168304 300012 168328
rect 297786 168272 299490 168304
rect 297725 168270 299490 168272
rect 97441 168267 97507 168270
rect 297725 168267 297791 168270
rect 99281 168058 99347 168061
rect 99422 168058 100004 168092
rect 99281 168056 100004 168058
rect 99281 168000 99286 168056
rect 99342 168032 100004 168056
rect 297633 168058 297699 168061
rect 299430 168058 300012 168092
rect 297633 168056 300012 168058
rect 99342 168000 99482 168032
rect 99281 167998 99482 168000
rect 297633 168000 297638 168056
rect 297694 168032 300012 168056
rect 297694 168000 299490 168032
rect 297633 167998 299490 168000
rect 99281 167995 99347 167998
rect 297633 167995 297699 167998
rect 291694 166228 291700 166292
rect 291764 166290 291770 166292
rect 292389 166290 292455 166293
rect 291764 166288 292455 166290
rect 291764 166232 292394 166288
rect 292450 166232 292455 166288
rect 291764 166230 292455 166232
rect 291764 166228 291770 166230
rect 292389 166227 292455 166230
rect 583520 165732 584960 165972
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 153653 159900 153719 159901
rect 156045 159900 156111 159901
rect 153584 159898 153590 159900
rect 153562 159838 153590 159898
rect 153584 159836 153590 159838
rect 153654 159896 153719 159900
rect 156032 159898 156038 159900
rect 153654 159840 153658 159896
rect 153714 159840 153719 159896
rect 153654 159836 153719 159840
rect 155954 159838 156038 159898
rect 156102 159896 156111 159900
rect 156106 159840 156111 159896
rect 156032 159836 156038 159838
rect 156102 159836 156111 159840
rect 153653 159835 153719 159836
rect 156045 159835 156111 159836
rect 160921 159900 160987 159901
rect 175917 159900 175983 159901
rect 160921 159896 160934 159900
rect 160998 159898 161004 159900
rect 175888 159898 175894 159900
rect 160921 159840 160926 159896
rect 160921 159836 160934 159840
rect 160998 159838 161078 159898
rect 175826 159838 175894 159898
rect 175958 159896 175983 159900
rect 175978 159840 175983 159896
rect 160998 159836 161004 159838
rect 175888 159836 175894 159838
rect 175958 159836 175983 159840
rect 160921 159835 160987 159836
rect 175917 159835 175983 159836
rect 348233 159900 348299 159901
rect 350993 159900 351059 159901
rect 356053 159900 356119 159901
rect 348233 159896 348286 159900
rect 348350 159898 348356 159900
rect 348233 159840 348238 159896
rect 348233 159836 348286 159840
rect 348350 159838 348390 159898
rect 350993 159896 351006 159900
rect 351070 159898 351076 159900
rect 356032 159898 356038 159900
rect 350993 159840 350998 159896
rect 348350 159836 348356 159838
rect 350993 159836 351006 159840
rect 351070 159838 351150 159898
rect 355962 159838 356038 159898
rect 356102 159896 356119 159900
rect 356114 159840 356119 159896
rect 351070 159836 351076 159838
rect 356032 159836 356038 159838
rect 356102 159836 356119 159840
rect 348233 159835 348299 159836
rect 350993 159835 351059 159836
rect 356053 159835 356119 159836
rect 358445 159900 358511 159901
rect 360929 159900 360995 159901
rect 368289 159900 368355 159901
rect 358445 159896 358486 159900
rect 358550 159898 358556 159900
rect 358445 159840 358450 159896
rect 358445 159836 358486 159840
rect 358550 159838 358602 159898
rect 358550 159836 358556 159838
rect 360928 159836 360934 159900
rect 360998 159898 361004 159900
rect 368272 159898 368278 159900
rect 360998 159838 361086 159898
rect 368198 159838 368278 159898
rect 368342 159896 368355 159900
rect 368350 159840 368355 159896
rect 360998 159836 361004 159838
rect 368272 159836 368278 159838
rect 368342 159836 368355 159840
rect 358445 159835 358511 159836
rect 360929 159835 360995 159836
rect 368289 159835 368355 159836
rect 165981 159628 166047 159629
rect 165960 159626 165966 159628
rect 165890 159566 165966 159626
rect 166030 159624 166047 159628
rect 166042 159568 166047 159624
rect 165960 159564 165966 159566
rect 166030 159564 166047 159568
rect 165981 159563 166047 159564
rect 353569 159628 353635 159629
rect 365897 159628 365963 159629
rect 353569 159624 353590 159628
rect 353654 159626 353660 159628
rect 353569 159568 353574 159624
rect 353569 159564 353590 159568
rect 353654 159566 353726 159626
rect 365897 159624 365966 159628
rect 365897 159568 365902 159624
rect 365958 159568 365966 159624
rect 353654 159564 353660 159566
rect 365897 159564 365966 159568
rect 366030 159626 366036 159628
rect 366030 159566 366054 159626
rect 366030 159564 366036 159566
rect 353569 159563 353635 159564
rect 365897 159563 365963 159564
rect 200113 159354 200179 159357
rect 265617 159354 265683 159357
rect 200113 159352 265683 159354
rect 200113 159296 200118 159352
rect 200174 159296 265622 159352
rect 265678 159296 265683 159352
rect 200113 159294 265683 159296
rect 200113 159291 200179 159294
rect 265617 159291 265683 159294
rect 298277 159354 298343 159357
rect 373993 159354 374059 159357
rect 298277 159352 374059 159354
rect 298277 159296 298282 159352
rect 298338 159296 373998 159352
rect 374054 159296 374059 159352
rect 298277 159294 374059 159296
rect 298277 159291 298343 159294
rect 373993 159291 374059 159294
rect 128302 159156 128308 159220
rect 128372 159218 128378 159220
rect 238201 159218 238267 159221
rect 128372 159216 238267 159218
rect 128372 159160 238206 159216
rect 238262 159160 238267 159216
rect 128372 159158 238267 159160
rect 128372 159156 128378 159158
rect 238201 159155 238267 159158
rect 173382 159020 173388 159084
rect 173452 159082 173458 159084
rect 284702 159082 284708 159084
rect 173452 159022 284708 159082
rect 173452 159020 173458 159022
rect 284702 159020 284708 159022
rect 284772 159020 284778 159084
rect 163630 158884 163636 158948
rect 163700 158946 163706 158948
rect 282126 158946 282132 158948
rect 163700 158886 282132 158946
rect 163700 158884 163706 158886
rect 282126 158884 282132 158886
rect 282196 158884 282202 158948
rect 293350 158884 293356 158948
rect 293420 158946 293426 158948
rect 293861 158946 293927 158949
rect 293420 158944 293927 158946
rect 293420 158888 293866 158944
rect 293922 158888 293927 158944
rect 293420 158886 293927 158888
rect 293420 158884 293426 158886
rect 293861 158883 293927 158886
rect 289261 158812 289327 158813
rect 158478 158748 158484 158812
rect 158548 158810 158554 158812
rect 283414 158810 283420 158812
rect 158548 158750 283420 158810
rect 158548 158748 158554 158750
rect 283414 158748 283420 158750
rect 283484 158748 283490 158812
rect 289261 158810 289308 158812
rect 289216 158808 289308 158810
rect 289216 158752 289266 158808
rect 289216 158750 289308 158752
rect 289261 158748 289308 158750
rect 289372 158748 289378 158812
rect 293166 158748 293172 158812
rect 293236 158810 293242 158812
rect 293493 158810 293559 158813
rect 293236 158808 293559 158810
rect 293236 158752 293498 158808
rect 293554 158752 293559 158808
rect 293236 158750 293559 158752
rect 293236 158748 293242 158750
rect 289261 158747 289327 158748
rect 293493 158747 293559 158750
rect 298686 158748 298692 158812
rect 298756 158810 298762 158812
rect 299013 158810 299079 158813
rect 298756 158808 299079 158810
rect 298756 158752 299018 158808
rect 299074 158752 299079 158808
rect 298756 158750 299079 158752
rect 298756 158748 298762 158750
rect 299013 158747 299079 158750
rect 116209 158676 116275 158677
rect 118233 158676 118299 158677
rect 116158 158674 116164 158676
rect 116118 158614 116164 158674
rect 116228 158672 116275 158676
rect 118182 158674 118188 158676
rect 116270 158616 116275 158672
rect 116158 158612 116164 158614
rect 116228 158612 116275 158616
rect 118142 158614 118188 158674
rect 118252 158672 118299 158676
rect 118294 158616 118299 158672
rect 118182 158612 118188 158614
rect 118252 158612 118299 158616
rect 119654 158612 119660 158676
rect 119724 158674 119730 158676
rect 119889 158674 119955 158677
rect 120625 158676 120691 158677
rect 121913 158676 121979 158677
rect 126513 158676 126579 158677
rect 127617 158676 127683 158677
rect 128721 158676 128787 158677
rect 120574 158674 120580 158676
rect 119724 158672 119955 158674
rect 119724 158616 119894 158672
rect 119950 158616 119955 158672
rect 119724 158614 119955 158616
rect 120534 158614 120580 158674
rect 120644 158672 120691 158676
rect 121862 158674 121868 158676
rect 120686 158616 120691 158672
rect 119724 158612 119730 158614
rect 116209 158611 116275 158612
rect 118233 158611 118299 158612
rect 119889 158611 119955 158614
rect 120574 158612 120580 158614
rect 120644 158612 120691 158616
rect 121822 158614 121868 158674
rect 121932 158672 121979 158676
rect 126462 158674 126468 158676
rect 121974 158616 121979 158672
rect 121862 158612 121868 158614
rect 121932 158612 121979 158616
rect 126422 158614 126468 158674
rect 126532 158672 126579 158676
rect 127566 158674 127572 158676
rect 126574 158616 126579 158672
rect 126462 158612 126468 158614
rect 126532 158612 126579 158616
rect 127526 158614 127572 158674
rect 127636 158672 127683 158676
rect 128670 158674 128676 158676
rect 127678 158616 127683 158672
rect 127566 158612 127572 158614
rect 127636 158612 127683 158616
rect 128630 158614 128676 158674
rect 128740 158672 128787 158676
rect 128782 158616 128787 158672
rect 128670 158612 128676 158614
rect 128740 158612 128787 158616
rect 130142 158612 130148 158676
rect 130212 158674 130218 158676
rect 130561 158674 130627 158677
rect 131297 158676 131363 158677
rect 132401 158676 132467 158677
rect 133505 158676 133571 158677
rect 131246 158674 131252 158676
rect 130212 158672 130627 158674
rect 130212 158616 130566 158672
rect 130622 158616 130627 158672
rect 130212 158614 130627 158616
rect 131206 158614 131252 158674
rect 131316 158672 131363 158676
rect 132350 158674 132356 158676
rect 131358 158616 131363 158672
rect 130212 158612 130218 158614
rect 120625 158611 120691 158612
rect 121913 158611 121979 158612
rect 126513 158611 126579 158612
rect 127617 158611 127683 158612
rect 128721 158611 128787 158612
rect 130561 158611 130627 158614
rect 131246 158612 131252 158614
rect 131316 158612 131363 158616
rect 132310 158614 132356 158674
rect 132420 158672 132467 158676
rect 133454 158674 133460 158676
rect 132462 158616 132467 158672
rect 132350 158612 132356 158614
rect 132420 158612 132467 158616
rect 133414 158614 133460 158674
rect 133524 158672 133571 158676
rect 133566 158616 133571 158672
rect 133454 158612 133460 158614
rect 133524 158612 133571 158616
rect 138606 158612 138612 158676
rect 138676 158674 138682 158676
rect 139301 158674 139367 158677
rect 138676 158672 139367 158674
rect 138676 158616 139306 158672
rect 139362 158616 139367 158672
rect 138676 158614 139367 158616
rect 138676 158612 138682 158614
rect 131297 158611 131363 158612
rect 132401 158611 132467 158612
rect 133505 158611 133571 158612
rect 139301 158611 139367 158614
rect 159214 158612 159220 158676
rect 159284 158674 159290 158676
rect 159633 158674 159699 158677
rect 168281 158676 168347 158677
rect 188705 158676 188771 158677
rect 206001 158676 206067 158677
rect 168230 158674 168236 158676
rect 159284 158672 159699 158674
rect 159284 158616 159638 158672
rect 159694 158616 159699 158672
rect 159284 158614 159699 158616
rect 168190 158614 168236 158674
rect 168300 158672 168347 158676
rect 188654 158674 188660 158676
rect 168342 158616 168347 158672
rect 159284 158612 159290 158614
rect 159633 158611 159699 158614
rect 168230 158612 168236 158614
rect 168300 158612 168347 158616
rect 188614 158614 188660 158674
rect 188724 158672 188771 158676
rect 205950 158674 205956 158676
rect 188766 158616 188771 158672
rect 188654 158612 188660 158614
rect 188724 158612 188771 158616
rect 205910 158614 205956 158674
rect 206020 158672 206067 158676
rect 206062 158616 206067 158672
rect 205950 158612 205956 158614
rect 206020 158612 206067 158616
rect 315798 158612 315804 158676
rect 315868 158674 315874 158676
rect 316033 158674 316099 158677
rect 315868 158672 316099 158674
rect 315868 158616 316038 158672
rect 316094 158616 316099 158672
rect 315868 158614 316099 158616
rect 315868 158612 315874 158614
rect 168281 158611 168347 158612
rect 188705 158611 188771 158612
rect 206001 158611 206067 158612
rect 316033 158611 316099 158614
rect 317045 158676 317111 158677
rect 319437 158676 319503 158677
rect 320541 158676 320607 158677
rect 321645 158676 321711 158677
rect 323117 158676 323183 158677
rect 327533 158676 327599 158677
rect 328269 158676 328335 158677
rect 329925 158676 329991 158677
rect 317045 158672 317092 158676
rect 317156 158674 317162 158676
rect 317045 158616 317050 158672
rect 317045 158612 317092 158616
rect 317156 158614 317202 158674
rect 319437 158672 319484 158676
rect 319548 158674 319554 158676
rect 319437 158616 319442 158672
rect 317156 158612 317162 158614
rect 319437 158612 319484 158616
rect 319548 158614 319594 158674
rect 320541 158672 320588 158676
rect 320652 158674 320658 158676
rect 320541 158616 320546 158672
rect 319548 158612 319554 158614
rect 320541 158612 320588 158616
rect 320652 158614 320698 158674
rect 321645 158672 321692 158676
rect 321756 158674 321762 158676
rect 321645 158616 321650 158672
rect 320652 158612 320658 158614
rect 321645 158612 321692 158616
rect 321756 158614 321802 158674
rect 323117 158672 323164 158676
rect 323228 158674 323234 158676
rect 323117 158616 323122 158672
rect 321756 158612 321762 158614
rect 323117 158612 323164 158616
rect 323228 158614 323274 158674
rect 327533 158672 327580 158676
rect 327644 158674 327650 158676
rect 327533 158616 327538 158672
rect 323228 158612 323234 158614
rect 327533 158612 327580 158616
rect 327644 158614 327690 158674
rect 328269 158672 328316 158676
rect 328380 158674 328386 158676
rect 328269 158616 328274 158672
rect 327644 158612 327650 158614
rect 328269 158612 328316 158616
rect 328380 158614 328426 158674
rect 329925 158672 329972 158676
rect 330036 158674 330042 158676
rect 330293 158674 330359 158677
rect 331213 158676 331279 158677
rect 332317 158676 332383 158677
rect 333605 158676 333671 158677
rect 334525 158676 334591 158677
rect 335813 158676 335879 158677
rect 335997 158676 336063 158677
rect 336917 158676 336983 158677
rect 338389 158676 338455 158677
rect 339309 158676 339375 158677
rect 340965 158676 341031 158677
rect 343541 158676 343607 158677
rect 347589 158676 347655 158677
rect 354397 158676 354463 158677
rect 330702 158674 330708 158676
rect 329925 158616 329930 158672
rect 328380 158612 328386 158614
rect 329925 158612 329972 158616
rect 330036 158614 330082 158674
rect 330293 158672 330708 158674
rect 330293 158616 330298 158672
rect 330354 158616 330708 158672
rect 330293 158614 330708 158616
rect 330036 158612 330042 158614
rect 317045 158611 317111 158612
rect 319437 158611 319503 158612
rect 320541 158611 320607 158612
rect 321645 158611 321711 158612
rect 323117 158611 323183 158612
rect 327533 158611 327599 158612
rect 328269 158611 328335 158612
rect 329925 158611 329991 158612
rect 330293 158611 330359 158614
rect 330702 158612 330708 158614
rect 330772 158612 330778 158676
rect 331213 158672 331260 158676
rect 331324 158674 331330 158676
rect 331213 158616 331218 158672
rect 331213 158612 331260 158616
rect 331324 158614 331370 158674
rect 332317 158672 332364 158676
rect 332428 158674 332434 158676
rect 332317 158616 332322 158672
rect 331324 158612 331330 158614
rect 332317 158612 332364 158616
rect 332428 158614 332474 158674
rect 333605 158672 333652 158676
rect 333716 158674 333722 158676
rect 333605 158616 333610 158672
rect 332428 158612 332434 158614
rect 333605 158612 333652 158616
rect 333716 158614 333762 158674
rect 334525 158672 334572 158676
rect 334636 158674 334642 158676
rect 335813 158674 335860 158676
rect 334525 158616 334530 158672
rect 333716 158612 333722 158614
rect 334525 158612 334572 158616
rect 334636 158614 334682 158674
rect 335768 158672 335860 158674
rect 335768 158616 335818 158672
rect 335768 158614 335860 158616
rect 334636 158612 334642 158614
rect 335813 158612 335860 158614
rect 335924 158612 335930 158676
rect 335997 158672 336044 158676
rect 336108 158674 336114 158676
rect 335997 158616 336002 158672
rect 335997 158612 336044 158616
rect 336108 158614 336154 158674
rect 336917 158672 336964 158676
rect 337028 158674 337034 158676
rect 336917 158616 336922 158672
rect 336108 158612 336114 158614
rect 336917 158612 336964 158616
rect 337028 158614 337074 158674
rect 338389 158672 338436 158676
rect 338500 158674 338506 158676
rect 338389 158616 338394 158672
rect 337028 158612 337034 158614
rect 338389 158612 338436 158616
rect 338500 158614 338546 158674
rect 339309 158672 339356 158676
rect 339420 158674 339426 158676
rect 339309 158616 339314 158672
rect 338500 158612 338506 158614
rect 339309 158612 339356 158616
rect 339420 158614 339466 158674
rect 340965 158672 341012 158676
rect 341076 158674 341082 158676
rect 340965 158616 340970 158672
rect 339420 158612 339426 158614
rect 340965 158612 341012 158616
rect 341076 158614 341122 158674
rect 343541 158672 343588 158676
rect 343652 158674 343658 158676
rect 343541 158616 343546 158672
rect 341076 158612 341082 158614
rect 343541 158612 343588 158616
rect 343652 158614 343698 158674
rect 347589 158672 347636 158676
rect 347700 158674 347706 158676
rect 347589 158616 347594 158672
rect 343652 158612 343658 158614
rect 347589 158612 347636 158616
rect 347700 158614 347746 158674
rect 354397 158672 354444 158676
rect 354508 158674 354514 158676
rect 355225 158674 355291 158677
rect 356973 158676 357039 158677
rect 363413 158676 363479 158677
rect 370957 158676 371023 158677
rect 373441 158676 373507 158677
rect 376017 158676 376083 158677
rect 378593 158676 378659 158677
rect 380985 158676 381051 158677
rect 383561 158676 383627 158677
rect 385953 158676 386019 158677
rect 388529 158676 388595 158677
rect 355726 158674 355732 158676
rect 354397 158616 354402 158672
rect 347700 158612 347706 158614
rect 354397 158612 354444 158616
rect 354508 158614 354554 158674
rect 355225 158672 355732 158674
rect 355225 158616 355230 158672
rect 355286 158616 355732 158672
rect 355225 158614 355732 158616
rect 354508 158612 354514 158614
rect 331213 158611 331279 158612
rect 332317 158611 332383 158612
rect 333605 158611 333671 158612
rect 334525 158611 334591 158612
rect 335813 158611 335879 158612
rect 335997 158611 336063 158612
rect 336917 158611 336983 158612
rect 338389 158611 338455 158612
rect 339309 158611 339375 158612
rect 340965 158611 341031 158612
rect 343541 158611 343607 158612
rect 347589 158611 347655 158612
rect 354397 158611 354463 158612
rect 355225 158611 355291 158614
rect 355726 158612 355732 158614
rect 355796 158612 355802 158676
rect 356973 158672 357020 158676
rect 357084 158674 357090 158676
rect 356973 158616 356978 158672
rect 356973 158612 357020 158616
rect 357084 158614 357130 158674
rect 363413 158672 363460 158676
rect 363524 158674 363530 158676
rect 363413 158616 363418 158672
rect 357084 158612 357090 158614
rect 363413 158612 363460 158616
rect 363524 158614 363570 158674
rect 370957 158672 371004 158676
rect 371068 158674 371074 158676
rect 373390 158674 373396 158676
rect 370957 158616 370962 158672
rect 363524 158612 363530 158614
rect 370957 158612 371004 158616
rect 371068 158614 371114 158674
rect 373350 158614 373396 158674
rect 373460 158672 373507 158676
rect 375966 158674 375972 158676
rect 373502 158616 373507 158672
rect 371068 158612 371074 158614
rect 373390 158612 373396 158614
rect 373460 158612 373507 158616
rect 375926 158614 375972 158674
rect 376036 158672 376083 158676
rect 378542 158674 378548 158676
rect 376078 158616 376083 158672
rect 375966 158612 375972 158614
rect 376036 158612 376083 158616
rect 378502 158614 378548 158674
rect 378612 158672 378659 158676
rect 380934 158674 380940 158676
rect 378654 158616 378659 158672
rect 378542 158612 378548 158614
rect 378612 158612 378659 158616
rect 380894 158614 380940 158674
rect 381004 158672 381051 158676
rect 383510 158674 383516 158676
rect 381046 158616 381051 158672
rect 380934 158612 380940 158614
rect 381004 158612 381051 158616
rect 383470 158614 383516 158674
rect 383580 158672 383627 158676
rect 385902 158674 385908 158676
rect 383622 158616 383627 158672
rect 383510 158612 383516 158614
rect 383580 158612 383627 158616
rect 385862 158614 385908 158674
rect 385972 158672 386019 158676
rect 388478 158674 388484 158676
rect 386014 158616 386019 158672
rect 385902 158612 385908 158614
rect 385972 158612 386019 158616
rect 388438 158614 388484 158674
rect 388548 158672 388595 158676
rect 388590 158616 388595 158672
rect 388478 158612 388484 158614
rect 388548 158612 388595 158616
rect 391054 158612 391060 158676
rect 391124 158674 391130 158676
rect 391473 158674 391539 158677
rect 391124 158672 391539 158674
rect 391124 158616 391478 158672
rect 391534 158616 391539 158672
rect 391124 158614 391539 158616
rect 391124 158612 391130 158614
rect 356973 158611 357039 158612
rect 363413 158611 363479 158612
rect 370957 158611 371023 158612
rect 373441 158611 373507 158612
rect 376017 158611 376083 158612
rect 378593 158611 378659 158612
rect 380985 158611 381051 158612
rect 383561 158611 383627 158612
rect 385953 158611 386019 158612
rect 388529 158611 388595 158612
rect 391473 158611 391539 158614
rect 393446 158612 393452 158676
rect 393516 158674 393522 158676
rect 394233 158674 394299 158677
rect 395889 158676 395955 158677
rect 398465 158676 398531 158677
rect 401041 158676 401107 158677
rect 395838 158674 395844 158676
rect 393516 158672 394299 158674
rect 393516 158616 394238 158672
rect 394294 158616 394299 158672
rect 393516 158614 394299 158616
rect 395798 158614 395844 158674
rect 395908 158672 395955 158676
rect 398414 158674 398420 158676
rect 395950 158616 395955 158672
rect 393516 158612 393522 158614
rect 394233 158611 394299 158614
rect 395838 158612 395844 158614
rect 395908 158612 395955 158616
rect 398374 158614 398420 158674
rect 398484 158672 398531 158676
rect 400990 158674 400996 158676
rect 398526 158616 398531 158672
rect 398414 158612 398420 158614
rect 398484 158612 398531 158616
rect 400950 158614 400996 158674
rect 401060 158672 401107 158676
rect 401102 158616 401107 158672
rect 400990 158612 400996 158614
rect 401060 158612 401107 158616
rect 403382 158612 403388 158676
rect 403452 158674 403458 158676
rect 403985 158674 404051 158677
rect 403452 158672 404051 158674
rect 403452 158616 403990 158672
rect 404046 158616 404051 158672
rect 403452 158614 404051 158616
rect 403452 158612 403458 158614
rect 395889 158611 395955 158612
rect 398465 158611 398531 158612
rect 401041 158611 401107 158612
rect 403985 158611 404051 158614
rect 405958 158612 405964 158676
rect 406028 158674 406034 158676
rect 406469 158674 406535 158677
rect 406028 158672 406535 158674
rect 406028 158616 406474 158672
rect 406530 158616 406535 158672
rect 406028 158614 406535 158616
rect 406028 158612 406034 158614
rect 406469 158611 406535 158614
rect 135897 158540 135963 158541
rect 137001 158540 137067 158541
rect 135846 158538 135852 158540
rect 135806 158478 135852 158538
rect 135916 158536 135963 158540
rect 136950 158538 136956 158540
rect 135958 158480 135963 158536
rect 135846 158476 135852 158478
rect 135916 158476 135963 158480
rect 136910 158478 136956 158538
rect 137020 158536 137067 158540
rect 137062 158480 137067 158536
rect 136950 158476 136956 158478
rect 137020 158476 137067 158480
rect 138054 158476 138060 158540
rect 138124 158538 138130 158540
rect 138381 158538 138447 158541
rect 138124 158536 138447 158538
rect 138124 158480 138386 158536
rect 138442 158480 138447 158536
rect 138124 158478 138447 158480
rect 138124 158476 138130 158478
rect 135897 158475 135963 158476
rect 137001 158475 137067 158476
rect 138381 158475 138447 158478
rect 139526 158476 139532 158540
rect 139596 158538 139602 158540
rect 139669 158538 139735 158541
rect 139596 158536 139735 158538
rect 139596 158480 139674 158536
rect 139730 158480 139735 158536
rect 139596 158478 139735 158480
rect 139596 158476 139602 158478
rect 139669 158475 139735 158478
rect 158110 158476 158116 158540
rect 158180 158538 158186 158540
rect 278681 158538 278747 158541
rect 358118 158538 358124 158540
rect 158180 158536 358124 158538
rect 158180 158480 278686 158536
rect 278742 158480 358124 158536
rect 158180 158478 358124 158480
rect 158180 158476 158186 158478
rect 278681 158475 278747 158478
rect 358118 158476 358124 158478
rect 358188 158476 358194 158540
rect 183502 158340 183508 158404
rect 183572 158402 183578 158404
rect 184013 158402 184079 158405
rect 185945 158404 186011 158405
rect 185894 158402 185900 158404
rect 183572 158400 184079 158402
rect 183572 158344 184018 158400
rect 184074 158344 184079 158400
rect 183572 158342 184079 158344
rect 185854 158342 185900 158402
rect 185964 158400 186011 158404
rect 186006 158344 186011 158400
rect 183572 158340 183578 158342
rect 184013 158339 184079 158342
rect 185894 158340 185900 158342
rect 185964 158340 186011 158344
rect 193438 158340 193444 158404
rect 193508 158402 193514 158404
rect 276013 158402 276079 158405
rect 277117 158402 277183 158405
rect 328678 158402 328684 158404
rect 193508 158342 200130 158402
rect 193508 158340 193514 158342
rect 185945 158339 186011 158340
rect 123150 158204 123156 158268
rect 123220 158266 123226 158268
rect 123937 158266 124003 158269
rect 134609 158268 134675 158269
rect 134558 158266 134564 158268
rect 123220 158264 124003 158266
rect 123220 158208 123942 158264
rect 123998 158208 124003 158264
rect 123220 158206 124003 158208
rect 134518 158206 134564 158266
rect 134628 158264 134675 158268
rect 134670 158208 134675 158264
rect 123220 158204 123226 158206
rect 123937 158203 124003 158206
rect 134558 158204 134564 158206
rect 134628 158204 134675 158208
rect 141182 158204 141188 158268
rect 141252 158266 141258 158268
rect 141509 158266 141575 158269
rect 141785 158268 141851 158269
rect 146017 158268 146083 158269
rect 146385 158268 146451 158269
rect 150985 158268 151051 158269
rect 141734 158266 141740 158268
rect 141252 158264 141575 158266
rect 141252 158208 141514 158264
rect 141570 158208 141575 158264
rect 141252 158206 141575 158208
rect 141694 158206 141740 158266
rect 141804 158264 141851 158268
rect 145966 158266 145972 158268
rect 141846 158208 141851 158264
rect 141252 158204 141258 158206
rect 134609 158203 134675 158204
rect 141509 158203 141575 158206
rect 141734 158204 141740 158206
rect 141804 158204 141851 158208
rect 145926 158206 145972 158266
rect 146036 158264 146083 158268
rect 146334 158266 146340 158268
rect 146078 158208 146083 158264
rect 145966 158204 145972 158206
rect 146036 158204 146083 158208
rect 146294 158206 146340 158266
rect 146404 158264 146451 158268
rect 150934 158266 150940 158268
rect 146446 158208 146451 158264
rect 146334 158204 146340 158206
rect 146404 158204 146451 158208
rect 150894 158206 150940 158266
rect 151004 158264 151051 158268
rect 151046 158208 151051 158264
rect 150934 158204 150940 158206
rect 151004 158204 151051 158208
rect 191046 158204 191052 158268
rect 191116 158266 191122 158268
rect 191465 158266 191531 158269
rect 195881 158268 195947 158269
rect 195830 158266 195836 158268
rect 191116 158264 191531 158266
rect 191116 158208 191470 158264
rect 191526 158208 191531 158264
rect 191116 158206 191531 158208
rect 195790 158206 195836 158266
rect 195900 158264 195947 158268
rect 195942 158208 195947 158264
rect 191116 158204 191122 158206
rect 141785 158203 141851 158204
rect 146017 158203 146083 158204
rect 146385 158203 146451 158204
rect 150985 158203 151051 158204
rect 191465 158203 191531 158206
rect 195830 158204 195836 158206
rect 195900 158204 195947 158208
rect 200070 158266 200130 158342
rect 276013 158400 328684 158402
rect 276013 158344 276018 158400
rect 276074 158344 277122 158400
rect 277178 158344 328684 158400
rect 276013 158342 328684 158344
rect 276013 158339 276079 158342
rect 277117 158339 277183 158342
rect 328678 158340 328684 158342
rect 328748 158340 328754 158404
rect 278313 158266 278379 158269
rect 200070 158264 278379 158266
rect 200070 158208 278318 158264
rect 278374 158208 278379 158264
rect 200070 158206 278379 158208
rect 195881 158203 195947 158204
rect 278313 158203 278379 158206
rect 283833 158266 283899 158269
rect 338113 158268 338179 158269
rect 333462 158266 333468 158268
rect 283833 158264 333468 158266
rect 283833 158208 283838 158264
rect 283894 158208 333468 158264
rect 283833 158206 333468 158208
rect 283833 158203 283899 158206
rect 333462 158204 333468 158206
rect 333532 158204 333538 158268
rect 338062 158266 338068 158268
rect 338022 158206 338068 158266
rect 338132 158264 338179 158268
rect 338174 158208 338179 158264
rect 338062 158204 338068 158206
rect 338132 158204 338179 158208
rect 338113 158203 338179 158204
rect 343909 158268 343975 158269
rect 348693 158268 348759 158269
rect 353293 158268 353359 158269
rect 343909 158264 343956 158268
rect 344020 158266 344026 158268
rect 343909 158208 343914 158264
rect 343909 158204 343956 158208
rect 344020 158206 344066 158266
rect 348693 158264 348740 158268
rect 348804 158266 348810 158268
rect 348693 158208 348698 158264
rect 344020 158204 344026 158206
rect 348693 158204 348740 158208
rect 348804 158206 348850 158266
rect 353293 158264 353340 158268
rect 353404 158266 353410 158268
rect 353293 158208 353298 158264
rect 348804 158204 348810 158206
rect 353293 158204 353340 158208
rect 353404 158206 353450 158266
rect 353404 158204 353410 158206
rect 343909 158203 343975 158204
rect 348693 158203 348759 158204
rect 353293 158203 353359 158204
rect 117078 158068 117084 158132
rect 117148 158130 117154 158132
rect 117221 158130 117287 158133
rect 117148 158128 117287 158130
rect 117148 158072 117226 158128
rect 117282 158072 117287 158128
rect 117148 158070 117287 158072
rect 117148 158068 117154 158070
rect 117221 158067 117287 158070
rect 147622 158068 147628 158132
rect 147692 158130 147698 158132
rect 148685 158130 148751 158133
rect 147692 158128 148751 158130
rect 147692 158072 148690 158128
rect 148746 158072 148751 158128
rect 147692 158070 148751 158072
rect 147692 158068 147698 158070
rect 148685 158067 148751 158070
rect 170990 158068 170996 158132
rect 171060 158130 171066 158132
rect 238293 158130 238359 158133
rect 171060 158128 238359 158130
rect 171060 158072 238298 158128
rect 238354 158072 238359 158128
rect 171060 158070 238359 158072
rect 171060 158068 171066 158070
rect 238293 158067 238359 158070
rect 276565 158130 276631 158133
rect 326470 158130 326476 158132
rect 276565 158128 326476 158130
rect 276565 158072 276570 158128
rect 276626 158072 326476 158128
rect 276565 158070 326476 158072
rect 276565 158067 276631 158070
rect 326470 158068 326476 158070
rect 326540 158068 326546 158132
rect 140681 157996 140747 157997
rect 140630 157994 140636 157996
rect 140590 157934 140636 157994
rect 140700 157992 140747 157996
rect 140742 157936 140747 157992
rect 140630 157932 140636 157934
rect 140700 157932 140747 157936
rect 142838 157932 142844 157996
rect 142908 157994 142914 157996
rect 143073 157994 143139 157997
rect 142908 157992 143139 157994
rect 142908 157936 143078 157992
rect 143134 157936 143139 157992
rect 142908 157934 143139 157936
rect 142908 157932 142914 157934
rect 140681 157931 140747 157932
rect 143073 157931 143139 157934
rect 143574 157932 143580 157996
rect 143644 157994 143650 157996
rect 144545 157994 144611 157997
rect 143644 157992 144611 157994
rect 143644 157936 144550 157992
rect 144606 157936 144611 157992
rect 143644 157934 144611 157936
rect 143644 157932 143650 157934
rect 144545 157931 144611 157934
rect 290917 157994 290983 157997
rect 318190 157994 318196 157996
rect 290917 157992 318196 157994
rect 290917 157936 290922 157992
rect 290978 157936 318196 157992
rect 290917 157934 318196 157936
rect 290917 157931 290983 157934
rect 318190 157932 318196 157934
rect 318260 157932 318266 157996
rect 341149 157994 341215 157997
rect 341742 157994 341748 157996
rect 341149 157992 341748 157994
rect 341149 157936 341154 157992
rect 341210 157936 341748 157992
rect 341149 157934 341748 157936
rect 341149 157931 341215 157934
rect 341742 157932 341748 157934
rect 341812 157932 341818 157996
rect 345105 157994 345171 157997
rect 346393 157996 346459 157997
rect 345238 157994 345244 157996
rect 345105 157992 345244 157994
rect 345105 157936 345110 157992
rect 345166 157936 345244 157992
rect 345105 157934 345244 157936
rect 345105 157931 345171 157934
rect 345238 157932 345244 157934
rect 345308 157932 345314 157996
rect 346342 157994 346348 157996
rect 346302 157934 346348 157994
rect 346412 157992 346459 157996
rect 346454 157936 346459 157992
rect 346342 157932 346348 157934
rect 346412 157932 346459 157936
rect 346393 157931 346459 157932
rect 324221 157860 324287 157861
rect 130694 157796 130700 157860
rect 130764 157858 130770 157860
rect 283782 157858 283788 157860
rect 130764 157798 283788 157858
rect 130764 157796 130770 157798
rect 283782 157796 283788 157798
rect 283852 157796 283858 157860
rect 324221 157856 324268 157860
rect 324332 157858 324338 157860
rect 339585 157858 339651 157861
rect 340638 157858 340644 157860
rect 324221 157800 324226 157856
rect 324221 157796 324268 157800
rect 324332 157798 324378 157858
rect 339585 157856 340644 157858
rect 339585 157800 339590 157856
rect 339646 157800 340644 157856
rect 339585 157798 340644 157800
rect 324332 157796 324338 157798
rect 324221 157795 324287 157796
rect 339585 157795 339651 157798
rect 340638 157796 340644 157798
rect 340708 157796 340714 157860
rect 342345 157858 342411 157861
rect 342846 157858 342852 157860
rect 342345 157856 342852 157858
rect 342345 157800 342350 157856
rect 342406 157800 342852 157856
rect 342345 157798 342852 157800
rect 342345 157795 342411 157798
rect 342846 157796 342852 157798
rect 342916 157796 342922 157860
rect 145281 157724 145347 157725
rect 148409 157724 148475 157725
rect 148777 157724 148843 157725
rect 145230 157722 145236 157724
rect 145190 157662 145236 157722
rect 145300 157720 145347 157724
rect 148358 157722 148364 157724
rect 145342 157664 145347 157720
rect 145230 157660 145236 157662
rect 145300 157660 145347 157664
rect 148318 157662 148364 157722
rect 148428 157720 148475 157724
rect 148726 157722 148732 157724
rect 148470 157664 148475 157720
rect 148358 157660 148364 157662
rect 148428 157660 148475 157664
rect 148686 157662 148732 157722
rect 148796 157720 148843 157724
rect 148838 157664 148843 157720
rect 148726 157660 148732 157662
rect 148796 157660 148843 157664
rect 178534 157660 178540 157724
rect 178604 157722 178610 157724
rect 283598 157722 283604 157724
rect 178604 157662 283604 157722
rect 178604 157660 178610 157662
rect 283598 157660 283604 157662
rect 283668 157660 283674 157724
rect 145281 157659 145347 157660
rect 148409 157659 148475 157660
rect 148777 157659 148843 157660
rect 124254 157524 124260 157588
rect 124324 157586 124330 157588
rect 124765 157586 124831 157589
rect 155769 157588 155835 157589
rect 201033 157588 201099 157589
rect 203425 157588 203491 157589
rect 155718 157586 155724 157588
rect 124324 157584 124831 157586
rect 124324 157528 124770 157584
rect 124826 157528 124831 157584
rect 124324 157526 124831 157528
rect 155678 157526 155724 157586
rect 155788 157584 155835 157588
rect 200982 157586 200988 157588
rect 155830 157528 155835 157584
rect 124324 157524 124330 157526
rect 124765 157523 124831 157526
rect 155718 157524 155724 157526
rect 155788 157524 155835 157528
rect 200942 157526 200988 157586
rect 201052 157584 201099 157588
rect 203374 157586 203380 157588
rect 201094 157528 201099 157584
rect 200982 157524 200988 157526
rect 201052 157524 201099 157528
rect 203334 157526 203380 157586
rect 203444 157584 203491 157588
rect 203486 157528 203491 157584
rect 203374 157524 203380 157526
rect 203444 157524 203491 157528
rect 155769 157523 155835 157524
rect 201033 157523 201099 157524
rect 203425 157523 203491 157524
rect 285121 157586 285187 157589
rect 359222 157586 359228 157588
rect 285121 157584 359228 157586
rect 285121 157528 285126 157584
rect 285182 157528 359228 157584
rect 285121 157526 359228 157528
rect 285121 157523 285187 157526
rect 359222 157524 359228 157526
rect 359292 157524 359298 157588
rect 125409 157452 125475 157453
rect 133689 157452 133755 157453
rect 136081 157452 136147 157453
rect 143993 157452 144059 157453
rect 149881 157452 149947 157453
rect 151353 157452 151419 157453
rect 125358 157450 125364 157452
rect 125318 157390 125364 157450
rect 125428 157448 125475 157452
rect 133638 157450 133644 157452
rect 125470 157392 125475 157448
rect 125358 157388 125364 157390
rect 125428 157388 125475 157392
rect 133598 157390 133644 157450
rect 133708 157448 133755 157452
rect 136030 157450 136036 157452
rect 133750 157392 133755 157448
rect 133638 157388 133644 157390
rect 133708 157388 133755 157392
rect 135990 157390 136036 157450
rect 136100 157448 136147 157452
rect 143942 157450 143948 157452
rect 136142 157392 136147 157448
rect 136030 157388 136036 157390
rect 136100 157388 136147 157392
rect 143902 157390 143948 157450
rect 144012 157448 144059 157452
rect 149830 157450 149836 157452
rect 144054 157392 144059 157448
rect 143942 157388 143948 157390
rect 144012 157388 144059 157392
rect 149790 157390 149836 157450
rect 149900 157448 149947 157452
rect 151302 157450 151308 157452
rect 149942 157392 149947 157448
rect 149830 157388 149836 157390
rect 149900 157388 149947 157392
rect 151262 157390 151308 157450
rect 151372 157448 151419 157452
rect 151414 157392 151419 157448
rect 151302 157388 151308 157390
rect 151372 157388 151419 157392
rect 152222 157388 152228 157452
rect 152292 157450 152298 157452
rect 152641 157450 152707 157453
rect 152292 157448 152707 157450
rect 152292 157392 152646 157448
rect 152702 157392 152707 157448
rect 152292 157390 152707 157392
rect 152292 157388 152298 157390
rect 125409 157387 125475 157388
rect 133689 157387 133755 157388
rect 136081 157387 136147 157388
rect 143993 157387 144059 157388
rect 149881 157387 149947 157388
rect 151353 157387 151419 157388
rect 152641 157387 152707 157390
rect 153326 157388 153332 157452
rect 153396 157450 153402 157452
rect 153837 157450 153903 157453
rect 154481 157452 154547 157453
rect 157057 157452 157123 157453
rect 198457 157452 198523 157453
rect 295057 157452 295123 157453
rect 154430 157450 154436 157452
rect 153396 157448 153903 157450
rect 153396 157392 153842 157448
rect 153898 157392 153903 157448
rect 153396 157390 153903 157392
rect 154390 157390 154436 157450
rect 154500 157448 154547 157452
rect 157006 157450 157012 157452
rect 154542 157392 154547 157448
rect 153396 157388 153402 157390
rect 153837 157387 153903 157390
rect 154430 157388 154436 157390
rect 154500 157388 154547 157392
rect 156966 157390 157012 157450
rect 157076 157448 157123 157452
rect 157118 157392 157123 157448
rect 157006 157388 157012 157390
rect 157076 157388 157123 157392
rect 180926 157388 180932 157452
rect 180996 157388 181002 157452
rect 198406 157450 198412 157452
rect 198366 157390 198412 157450
rect 198476 157448 198523 157452
rect 295006 157450 295012 157452
rect 198518 157392 198523 157448
rect 198406 157388 198412 157390
rect 198476 157388 198523 157392
rect 294966 157390 295012 157450
rect 295076 157448 295123 157452
rect 295118 157392 295123 157448
rect 295006 157388 295012 157390
rect 295076 157388 295123 157392
rect 154481 157387 154547 157388
rect 157057 157387 157123 157388
rect 180934 157314 180994 157388
rect 198457 157387 198523 157388
rect 295057 157387 295123 157388
rect 324865 157450 324931 157453
rect 325366 157450 325372 157452
rect 324865 157448 325372 157450
rect 324865 157392 324870 157448
rect 324926 157392 325372 157448
rect 324865 157390 325372 157392
rect 324865 157387 324931 157390
rect 325366 157388 325372 157390
rect 325436 157388 325442 157452
rect 345749 157450 345815 157453
rect 349797 157452 349863 157453
rect 351085 157452 351151 157453
rect 352189 157452 352255 157453
rect 345974 157450 345980 157452
rect 345749 157448 345980 157450
rect 345749 157392 345754 157448
rect 345810 157392 345980 157448
rect 345749 157390 345980 157392
rect 345749 157387 345815 157390
rect 345974 157388 345980 157390
rect 346044 157388 346050 157452
rect 349797 157448 349844 157452
rect 349908 157450 349914 157452
rect 349797 157392 349802 157448
rect 349797 157388 349844 157392
rect 349908 157390 349954 157450
rect 351085 157448 351132 157452
rect 351196 157450 351202 157452
rect 351085 157392 351090 157448
rect 349908 157388 349914 157390
rect 351085 157388 351132 157392
rect 351196 157390 351242 157450
rect 352189 157448 352236 157452
rect 352300 157450 352306 157452
rect 352189 157392 352194 157448
rect 351196 157388 351202 157390
rect 352189 157388 352236 157392
rect 352300 157390 352346 157450
rect 352300 157388 352306 157390
rect 349797 157387 349863 157388
rect 351085 157387 351151 157388
rect 352189 157387 352255 157388
rect 281073 157314 281139 157317
rect 180934 157312 281139 157314
rect 180934 157256 281078 157312
rect 281134 157256 281139 157312
rect 180934 157254 281139 157256
rect 281073 157251 281139 157254
rect 207013 156906 207079 156909
rect 268193 156906 268259 156909
rect 207013 156904 268259 156906
rect 207013 156848 207018 156904
rect 207074 156848 268198 156904
rect 268254 156848 268259 156904
rect 207013 156846 268259 156848
rect 207013 156843 207079 156846
rect 268193 156843 268259 156846
rect 178033 156770 178099 156773
rect 260097 156770 260163 156773
rect 178033 156768 260163 156770
rect 178033 156712 178038 156768
rect 178094 156712 260102 156768
rect 260158 156712 260163 156768
rect 178033 156710 260163 156712
rect 178033 156707 178099 156710
rect 260097 156707 260163 156710
rect 290590 156708 290596 156772
rect 290660 156770 290666 156772
rect 290917 156770 290983 156773
rect 290660 156768 290983 156770
rect 290660 156712 290922 156768
rect 290978 156712 290983 156768
rect 290660 156710 290983 156712
rect 290660 156708 290666 156710
rect 290917 156707 290983 156710
rect 151813 156634 151879 156637
rect 258441 156634 258507 156637
rect 290733 156636 290799 156637
rect 290733 156634 290780 156636
rect 151813 156632 258507 156634
rect 151813 156576 151818 156632
rect 151874 156576 258446 156632
rect 258502 156576 258507 156632
rect 151813 156574 258507 156576
rect 290688 156632 290780 156634
rect 290688 156576 290738 156632
rect 290688 156574 290780 156576
rect 151813 156571 151879 156574
rect 258441 156571 258507 156574
rect 290733 156572 290780 156574
rect 290844 156572 290850 156636
rect 290733 156571 290799 156572
rect 139301 155954 139367 155957
rect 272609 155954 272675 155957
rect 139301 155952 272675 155954
rect 139301 155896 139306 155952
rect 139362 155896 272614 155952
rect 272670 155896 272675 155952
rect 139301 155894 272675 155896
rect 139301 155891 139367 155894
rect 272609 155891 272675 155894
rect 289486 155892 289492 155956
rect 289556 155954 289562 155956
rect 289629 155954 289695 155957
rect 289556 155952 289695 155954
rect 289556 155896 289634 155952
rect 289690 155896 289695 155952
rect 289556 155894 289695 155896
rect 289556 155892 289562 155894
rect 289629 155891 289695 155894
rect 144545 155818 144611 155821
rect 272793 155818 272859 155821
rect 144545 155816 272859 155818
rect 144545 155760 144550 155816
rect 144606 155760 272798 155816
rect 272854 155760 272859 155816
rect 144545 155758 272859 155760
rect 144545 155755 144611 155758
rect 272793 155755 272859 155758
rect 289118 155756 289124 155820
rect 289188 155818 289194 155820
rect 289445 155818 289511 155821
rect 289188 155816 289511 155818
rect 289188 155760 289450 155816
rect 289506 155760 289511 155816
rect 289188 155758 289511 155760
rect 289188 155756 289194 155758
rect 289445 155755 289511 155758
rect 224953 155546 225019 155549
rect 270953 155546 271019 155549
rect 224953 155544 271019 155546
rect 224953 155488 224958 155544
rect 225014 155488 270958 155544
rect 271014 155488 271019 155544
rect 224953 155486 271019 155488
rect 224953 155483 225019 155486
rect 270953 155483 271019 155486
rect 182173 155410 182239 155413
rect 262581 155410 262647 155413
rect 182173 155408 262647 155410
rect 182173 155352 182178 155408
rect 182234 155352 262586 155408
rect 262642 155352 262647 155408
rect 182173 155350 262647 155352
rect 182173 155347 182239 155350
rect 262581 155347 262647 155350
rect 160093 155274 160159 155277
rect 253381 155274 253447 155277
rect 160093 155272 253447 155274
rect 160093 155216 160098 155272
rect 160154 155216 253386 155272
rect 253442 155216 253447 155272
rect 160093 155214 253447 155216
rect 160093 155211 160159 155214
rect 253381 155211 253447 155214
rect 133689 154458 133755 154461
rect 275318 154458 275324 154460
rect 133689 154456 275324 154458
rect 133689 154400 133694 154456
rect 133750 154400 275324 154456
rect 133689 154398 275324 154400
rect 133689 154395 133755 154398
rect 275318 154396 275324 154398
rect 275388 154396 275394 154460
rect 136081 154322 136147 154325
rect 275134 154322 275140 154324
rect 136081 154320 275140 154322
rect 136081 154264 136086 154320
rect 136142 154264 275140 154320
rect 136081 154262 275140 154264
rect 136081 154259 136147 154262
rect 275134 154260 275140 154262
rect 275204 154260 275210 154324
rect 129733 153778 129799 153781
rect 254301 153778 254367 153781
rect 129733 153776 254367 153778
rect 129733 153720 129738 153776
rect 129794 153720 254306 153776
rect 254362 153720 254367 153776
rect 129733 153718 254367 153720
rect 129733 153715 129799 153718
rect 254301 153715 254367 153718
rect 288934 153036 288940 153100
rect 289004 153098 289010 153100
rect 289353 153098 289419 153101
rect 289004 153096 289419 153098
rect 289004 153040 289358 153096
rect 289414 153040 289419 153096
rect 289004 153038 289419 153040
rect 289004 153036 289010 153038
rect 289353 153035 289419 153038
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect 284886 152356 284892 152420
rect 284956 152418 284962 152420
rect 300853 152418 300919 152421
rect 284956 152416 300919 152418
rect 284956 152360 300858 152416
rect 300914 152360 300919 152416
rect 284956 152358 300919 152360
rect 284956 152356 284962 152358
rect 300853 152355 300919 152358
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 264329 148338 264395 148341
rect 277526 148338 277532 148340
rect 264329 148336 277532 148338
rect 264329 148280 264334 148336
rect 264390 148280 277532 148336
rect 264329 148278 277532 148280
rect 264329 148275 264395 148278
rect 277526 148276 277532 148278
rect 277596 148276 277602 148340
rect 273897 147658 273963 147661
rect 278998 147658 279004 147660
rect 273897 147656 279004 147658
rect 273897 147600 273902 147656
rect 273958 147600 279004 147656
rect 273897 147598 279004 147600
rect 273897 147595 273963 147598
rect 278998 147596 279004 147598
rect 279068 147596 279074 147660
rect 260097 141402 260163 141405
rect 277158 141402 277164 141404
rect 260097 141400 277164 141402
rect 260097 141344 260102 141400
rect 260158 141344 277164 141400
rect 260097 141342 277164 141344
rect 260097 141339 260163 141342
rect 277158 141340 277164 141342
rect 277228 141340 277234 141404
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 265157 129026 265223 129029
rect 278814 129026 278820 129028
rect 265157 129024 278820 129026
rect 265157 128968 265162 129024
rect 265218 128968 278820 129024
rect 265157 128966 278820 128968
rect 265157 128963 265223 128966
rect 278814 128964 278820 128966
rect 278884 128964 278890 129028
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 298318 80684 298324 80748
rect 298388 80746 298394 80748
rect 375373 80746 375439 80749
rect 298388 80744 375439 80746
rect 298388 80688 375378 80744
rect 375434 80688 375439 80744
rect 298388 80686 375439 80688
rect 298388 80684 298394 80686
rect 375373 80683 375439 80686
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 296478 18532 296484 18596
rect 296548 18594 296554 18596
rect 361573 18594 361639 18597
rect 296548 18592 361639 18594
rect 296548 18536 361578 18592
rect 361634 18536 361639 18592
rect 296548 18534 361639 18536
rect 296548 18532 296554 18534
rect 361573 18531 361639 18534
rect 287646 9556 287652 9620
rect 287716 9618 287722 9620
rect 383561 9618 383627 9621
rect 287716 9616 383627 9618
rect 287716 9560 383566 9616
rect 383622 9560 383627 9616
rect 287716 9558 383627 9560
rect 287716 9556 287722 9558
rect 383561 9555 383627 9558
rect 286542 9420 286548 9484
rect 286612 9482 286618 9484
rect 390645 9482 390711 9485
rect 286612 9480 390711 9482
rect 286612 9424 390650 9480
rect 390706 9424 390711 9480
rect 286612 9422 390711 9424
rect 286612 9420 286618 9422
rect 390645 9419 390711 9422
rect 286726 9284 286732 9348
rect 286796 9346 286802 9348
rect 404813 9346 404879 9349
rect 286796 9344 404879 9346
rect 286796 9288 404818 9344
rect 404874 9288 404879 9344
rect 286796 9286 404879 9288
rect 286796 9284 286802 9286
rect 404813 9283 404879 9286
rect 292246 9148 292252 9212
rect 292316 9210 292322 9212
rect 411897 9210 411963 9213
rect 292316 9208 411963 9210
rect 292316 9152 411902 9208
rect 411958 9152 411963 9208
rect 292316 9150 411963 9152
rect 292316 9148 292322 9150
rect 411897 9147 411963 9150
rect 288014 9012 288020 9076
rect 288084 9074 288090 9076
rect 408401 9074 408467 9077
rect 288084 9072 408467 9074
rect 288084 9016 408406 9072
rect 408462 9016 408467 9072
rect 288084 9014 408467 9016
rect 288084 9012 288090 9014
rect 408401 9011 408467 9014
rect 287830 8876 287836 8940
rect 287900 8938 287906 8940
rect 414289 8938 414355 8941
rect 287900 8936 414355 8938
rect 287900 8880 414294 8936
rect 414350 8880 414355 8936
rect 287900 8878 414355 8880
rect 287900 8876 287906 8878
rect 414289 8875 414355 8878
rect 293534 8740 293540 8804
rect 293604 8802 293610 8804
rect 387149 8802 387215 8805
rect 293604 8800 387215 8802
rect 293604 8744 387154 8800
rect 387210 8744 387215 8800
rect 293604 8742 387215 8744
rect 293604 8740 293610 8742
rect 387149 8739 387215 8742
rect 297398 6836 297404 6900
rect 297468 6898 297474 6900
rect 369393 6898 369459 6901
rect 297468 6896 369459 6898
rect 297468 6840 369398 6896
rect 369454 6840 369459 6896
rect 297468 6838 369459 6840
rect 297468 6836 297474 6838
rect 369393 6835 369459 6838
rect 298502 6700 298508 6764
rect 298572 6762 298578 6764
rect 375281 6762 375347 6765
rect 298572 6760 375347 6762
rect 298572 6704 375286 6760
rect 375342 6704 375347 6760
rect 298572 6702 375347 6704
rect 298572 6700 298578 6702
rect 375281 6699 375347 6702
rect -960 6490 480 6580
rect 282494 6564 282500 6628
rect 282564 6626 282570 6628
rect 367001 6626 367067 6629
rect 282564 6624 367067 6626
rect 282564 6568 367006 6624
rect 367062 6568 367067 6624
rect 282564 6566 367067 6568
rect 282564 6564 282570 6566
rect 367001 6563 367067 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 282678 6428 282684 6492
rect 282748 6490 282754 6492
rect 370589 6490 370655 6493
rect 282748 6488 370655 6490
rect 282748 6432 370594 6488
rect 370650 6432 370655 6488
rect 583520 6476 584960 6716
rect 282748 6430 370655 6432
rect 282748 6428 282754 6430
rect 370589 6427 370655 6430
rect 295926 6292 295932 6356
rect 295996 6354 296002 6356
rect 393037 6354 393103 6357
rect 295996 6352 393103 6354
rect 295996 6296 393042 6352
rect 393098 6296 393103 6352
rect 295996 6294 393103 6296
rect 295996 6292 296002 6294
rect 393037 6291 393103 6294
rect 292430 6156 292436 6220
rect 292500 6218 292506 6220
rect 389449 6218 389515 6221
rect 292500 6216 389515 6218
rect 292500 6160 389454 6216
rect 389510 6160 389515 6216
rect 292500 6158 389515 6160
rect 292500 6156 292506 6158
rect 389449 6155 389515 6158
rect 297582 6020 297588 6084
rect 297652 6082 297658 6084
rect 365805 6082 365871 6085
rect 297652 6080 365871 6082
rect 297652 6024 365810 6080
rect 365866 6024 365871 6080
rect 297652 6022 365871 6024
rect 297652 6020 297658 6022
rect 365805 6019 365871 6022
rect 297950 4932 297956 4996
rect 298020 4994 298026 4996
rect 364609 4994 364675 4997
rect 298020 4992 364675 4994
rect 298020 4936 364614 4992
rect 364670 4936 364675 4992
rect 298020 4934 364675 4936
rect 298020 4932 298026 4934
rect 364609 4931 364675 4934
rect 297766 4796 297772 4860
rect 297836 4858 297842 4860
rect 368197 4858 368263 4861
rect 297836 4856 368263 4858
rect 297836 4800 368202 4856
rect 368258 4800 368263 4856
rect 297836 4798 368263 4800
rect 297836 4796 297842 4798
rect 368197 4795 368263 4798
rect 296294 3980 296300 4044
rect 296364 4042 296370 4044
rect 384757 4042 384823 4045
rect 296364 4040 384823 4042
rect 296364 3984 384762 4040
rect 384818 3984 384823 4040
rect 296364 3982 384823 3984
rect 296364 3980 296370 3982
rect 384757 3979 384823 3982
rect 439446 3980 439452 4044
rect 439516 4042 439522 4044
rect 443821 4042 443887 4045
rect 439516 4040 443887 4042
rect 439516 3984 443826 4040
rect 443882 3984 443887 4040
rect 439516 3982 443887 3984
rect 439516 3980 439522 3982
rect 443821 3979 443887 3982
rect 286910 3844 286916 3908
rect 286980 3906 286986 3908
rect 379973 3906 380039 3909
rect 286980 3904 380039 3906
rect 286980 3848 379978 3904
rect 380034 3848 380039 3904
rect 286980 3846 380039 3848
rect 286980 3844 286986 3846
rect 379973 3843 380039 3846
rect 296110 3708 296116 3772
rect 296180 3770 296186 3772
rect 391841 3770 391907 3773
rect 296180 3768 391907 3770
rect 296180 3712 391846 3768
rect 391902 3712 391907 3768
rect 296180 3710 391907 3712
rect 296180 3708 296186 3710
rect 391841 3707 391907 3710
rect 295190 3572 295196 3636
rect 295260 3634 295266 3636
rect 397729 3634 397795 3637
rect 295260 3632 397795 3634
rect 295260 3576 397734 3632
rect 397790 3576 397795 3632
rect 295260 3574 397795 3576
rect 295260 3572 295266 3574
rect 397729 3571 397795 3574
rect 432045 3634 432111 3637
rect 437790 3634 437796 3636
rect 432045 3632 437796 3634
rect 432045 3576 432050 3632
rect 432106 3576 437796 3632
rect 432045 3574 437796 3576
rect 432045 3571 432111 3574
rect 437790 3572 437796 3574
rect 437860 3572 437866 3636
rect 293718 3436 293724 3500
rect 293788 3498 293794 3500
rect 398925 3498 398991 3501
rect 293788 3496 398991 3498
rect 293788 3440 398930 3496
rect 398986 3440 398991 3496
rect 293788 3438 398991 3440
rect 293788 3436 293794 3438
rect 398925 3435 398991 3438
rect 437422 3436 437428 3500
rect 437492 3498 437498 3500
rect 437933 3498 437999 3501
rect 439129 3500 439195 3501
rect 437492 3496 437999 3498
rect 437492 3440 437938 3496
rect 437994 3440 437999 3496
rect 437492 3438 437999 3440
rect 437492 3436 437498 3438
rect 437933 3435 437999 3438
rect 439078 3436 439084 3500
rect 439148 3498 439195 3500
rect 439148 3496 439240 3498
rect 439190 3440 439240 3496
rect 439148 3438 439240 3440
rect 439148 3436 439195 3438
rect 439129 3435 439195 3436
rect 288198 3300 288204 3364
rect 288268 3362 288274 3364
rect 394233 3362 394299 3365
rect 288268 3360 394299 3362
rect 288268 3304 394238 3360
rect 394294 3304 394299 3360
rect 288268 3302 394299 3304
rect 288268 3300 288274 3302
rect 394233 3299 394299 3302
rect 429653 3362 429719 3365
rect 437606 3362 437612 3364
rect 429653 3360 437612 3362
rect 429653 3304 429658 3360
rect 429714 3304 437612 3360
rect 429653 3302 437612 3304
rect 429653 3299 429719 3302
rect 437606 3300 437612 3302
rect 437676 3300 437682 3364
rect 285070 3164 285076 3228
rect 285140 3226 285146 3228
rect 363505 3226 363571 3229
rect 285140 3224 363571 3226
rect 285140 3168 363510 3224
rect 363566 3168 363571 3224
rect 285140 3166 363571 3168
rect 285140 3164 285146 3166
rect 363505 3163 363571 3166
<< via3 >>
rect 250668 477260 250732 477324
rect 268332 477260 268396 477324
rect 258028 477048 258092 477052
rect 258028 476992 258078 477048
rect 258078 476992 258092 477048
rect 258028 476988 258092 476992
rect 270908 476988 270972 477052
rect 305868 476988 305932 477052
rect 308444 476988 308508 477052
rect 243124 476852 243188 476916
rect 248276 476852 248340 476916
rect 253612 476852 253676 476916
rect 256188 476852 256252 476916
rect 278452 476852 278516 476916
rect 303476 476852 303540 476916
rect 311020 476852 311084 476916
rect 323348 476852 323412 476916
rect 325924 476852 325988 476916
rect 239628 476716 239692 476780
rect 257108 476716 257172 476780
rect 263548 476776 263612 476780
rect 263548 476720 263598 476776
rect 263598 476720 263612 476776
rect 263548 476716 263612 476720
rect 258396 476580 258460 476644
rect 260972 476580 261036 476644
rect 276060 476640 276124 476644
rect 276060 476584 276074 476640
rect 276074 476584 276124 476640
rect 276060 476580 276124 476584
rect 245332 476444 245396 476508
rect 262812 476444 262876 476508
rect 265940 476444 266004 476508
rect 313412 476444 313476 476508
rect 315804 476444 315868 476508
rect 235948 476368 236012 476372
rect 235948 476312 235998 476368
rect 235998 476312 236012 476368
rect 235948 476308 236012 476312
rect 244228 476368 244292 476372
rect 244228 476312 244278 476368
rect 244278 476312 244292 476368
rect 244228 476308 244292 476312
rect 248644 476308 248708 476372
rect 252324 476308 252388 476372
rect 254532 476308 254596 476372
rect 260788 476308 260852 476372
rect 263916 476308 263980 476372
rect 267596 476368 267660 476372
rect 267596 476312 267610 476368
rect 267610 476312 267660 476368
rect 267596 476308 267660 476312
rect 273484 476308 273548 476372
rect 274404 476368 274468 476372
rect 274404 476312 274454 476368
rect 274454 476312 274468 476368
rect 274404 476308 274468 476312
rect 318380 476308 318444 476372
rect 320956 476308 321020 476372
rect 237052 476172 237116 476236
rect 238156 476172 238220 476236
rect 240548 476172 240612 476236
rect 241836 476172 241900 476236
rect 246436 476172 246500 476236
rect 247540 476172 247604 476236
rect 250116 476172 250180 476236
rect 251404 476172 251468 476236
rect 253428 476172 253492 476236
rect 255820 476172 255884 476236
rect 259500 476172 259564 476236
rect 261708 476172 261772 476236
rect 265388 476172 265452 476236
rect 266492 476172 266556 476236
rect 268700 476172 268764 476236
rect 269804 476172 269868 476236
rect 271276 476172 271340 476236
rect 272196 476172 272260 476236
rect 273300 476172 273364 476236
rect 275876 476232 275940 476236
rect 275876 476176 275926 476232
rect 275926 476176 275940 476232
rect 275876 476172 275940 476176
rect 276980 476172 277044 476236
rect 278084 476172 278148 476236
rect 279188 476172 279252 476236
rect 280844 476172 280908 476236
rect 283420 476172 283484 476236
rect 285996 476172 286060 476236
rect 288204 476172 288268 476236
rect 290964 476172 291028 476236
rect 293356 476172 293420 476236
rect 295932 476172 295996 476236
rect 298508 476172 298572 476236
rect 300900 476232 300964 476236
rect 300900 476176 300950 476232
rect 300950 476176 300964 476232
rect 300900 476172 300964 476176
rect 282684 309028 282748 309092
rect 283420 308892 283484 308956
rect 282132 308756 282196 308820
rect 284708 308484 284772 308548
rect 297956 308212 298020 308276
rect 297404 308076 297468 308140
rect 277348 307940 277412 308004
rect 297588 307940 297652 308004
rect 298324 307940 298388 308004
rect 277532 307804 277596 307868
rect 278820 307864 278884 307868
rect 278820 307808 278834 307864
rect 278834 307808 278884 307864
rect 278820 307804 278884 307808
rect 279004 307804 279068 307868
rect 284892 307804 284956 307868
rect 296484 307804 296548 307868
rect 297772 307804 297836 307868
rect 298508 307804 298572 307868
rect 283788 306172 283852 306236
rect 283604 306036 283668 306100
rect 275324 303316 275388 303380
rect 275140 303180 275204 303244
rect 439452 302908 439516 302972
rect 439084 298692 439148 298756
rect 437428 287676 437492 287740
rect 287652 248100 287716 248164
rect 286916 247964 286980 248028
rect 289492 247828 289556 247892
rect 288204 247692 288268 247756
rect 286548 247556 286612 247620
rect 437612 247556 437676 247620
rect 295196 247420 295260 247484
rect 293540 247284 293604 247348
rect 286732 247072 286796 247076
rect 286732 247016 286782 247072
rect 286782 247016 286796 247072
rect 286732 247012 286796 247016
rect 287836 247072 287900 247076
rect 287836 247016 287886 247072
rect 287886 247016 287900 247072
rect 287836 247012 287900 247016
rect 288020 247072 288084 247076
rect 288020 247016 288070 247072
rect 288070 247016 288084 247072
rect 288020 247012 288084 247016
rect 288940 247072 289004 247076
rect 288940 247016 288990 247072
rect 288990 247016 289004 247072
rect 288940 247012 289004 247016
rect 289124 247072 289188 247076
rect 289124 247016 289174 247072
rect 289174 247016 289188 247072
rect 289124 247012 289188 247016
rect 290596 247072 290660 247076
rect 290596 247016 290646 247072
rect 290646 247016 290660 247072
rect 290596 247012 290660 247016
rect 292252 247012 292316 247076
rect 285076 246196 285140 246260
rect 295932 245380 295996 245444
rect 292436 245244 292500 245308
rect 437796 245244 437860 245308
rect 290780 245108 290844 245172
rect 293724 245108 293788 245172
rect 289308 244972 289372 245036
rect 282500 244836 282564 244900
rect 295012 244700 295076 244764
rect 296116 244700 296180 244764
rect 296300 244564 296364 244628
rect 293172 244428 293236 244492
rect 291700 244352 291764 244356
rect 291700 244296 291750 244352
rect 291750 244296 291764 244352
rect 291700 244292 291764 244296
rect 291884 244292 291948 244356
rect 293356 244292 293420 244356
rect 298140 244292 298204 244356
rect 298692 244352 298756 244356
rect 298692 244296 298742 244352
rect 298742 244296 298756 244352
rect 298692 244292 298756 244296
rect 291884 196012 291948 196076
rect 298140 187716 298204 187780
rect 291700 166228 291764 166292
rect 153590 159836 153654 159900
rect 156038 159896 156102 159900
rect 156038 159840 156050 159896
rect 156050 159840 156102 159896
rect 156038 159836 156102 159840
rect 160934 159896 160998 159900
rect 160934 159840 160982 159896
rect 160982 159840 160998 159896
rect 160934 159836 160998 159840
rect 175894 159896 175958 159900
rect 175894 159840 175922 159896
rect 175922 159840 175958 159896
rect 175894 159836 175958 159840
rect 348286 159896 348350 159900
rect 348286 159840 348294 159896
rect 348294 159840 348350 159896
rect 348286 159836 348350 159840
rect 351006 159896 351070 159900
rect 351006 159840 351054 159896
rect 351054 159840 351070 159896
rect 351006 159836 351070 159840
rect 356038 159896 356102 159900
rect 356038 159840 356058 159896
rect 356058 159840 356102 159896
rect 356038 159836 356102 159840
rect 358486 159896 358550 159900
rect 358486 159840 358506 159896
rect 358506 159840 358550 159896
rect 358486 159836 358550 159840
rect 360934 159896 360998 159900
rect 360934 159840 360990 159896
rect 360990 159840 360998 159896
rect 360934 159836 360998 159840
rect 368278 159896 368342 159900
rect 368278 159840 368294 159896
rect 368294 159840 368342 159896
rect 368278 159836 368342 159840
rect 165966 159624 166030 159628
rect 165966 159568 165986 159624
rect 165986 159568 166030 159624
rect 165966 159564 166030 159568
rect 353590 159624 353654 159628
rect 353590 159568 353630 159624
rect 353630 159568 353654 159624
rect 353590 159564 353654 159568
rect 365966 159564 366030 159628
rect 128308 159156 128372 159220
rect 173388 159020 173452 159084
rect 284708 159020 284772 159084
rect 163636 158884 163700 158948
rect 282132 158884 282196 158948
rect 293356 158884 293420 158948
rect 158484 158748 158548 158812
rect 283420 158748 283484 158812
rect 289308 158808 289372 158812
rect 289308 158752 289322 158808
rect 289322 158752 289372 158808
rect 289308 158748 289372 158752
rect 293172 158748 293236 158812
rect 298692 158748 298756 158812
rect 116164 158672 116228 158676
rect 116164 158616 116214 158672
rect 116214 158616 116228 158672
rect 116164 158612 116228 158616
rect 118188 158672 118252 158676
rect 118188 158616 118238 158672
rect 118238 158616 118252 158672
rect 118188 158612 118252 158616
rect 119660 158612 119724 158676
rect 120580 158672 120644 158676
rect 120580 158616 120630 158672
rect 120630 158616 120644 158672
rect 120580 158612 120644 158616
rect 121868 158672 121932 158676
rect 121868 158616 121918 158672
rect 121918 158616 121932 158672
rect 121868 158612 121932 158616
rect 126468 158672 126532 158676
rect 126468 158616 126518 158672
rect 126518 158616 126532 158672
rect 126468 158612 126532 158616
rect 127572 158672 127636 158676
rect 127572 158616 127622 158672
rect 127622 158616 127636 158672
rect 127572 158612 127636 158616
rect 128676 158672 128740 158676
rect 128676 158616 128726 158672
rect 128726 158616 128740 158672
rect 128676 158612 128740 158616
rect 130148 158612 130212 158676
rect 131252 158672 131316 158676
rect 131252 158616 131302 158672
rect 131302 158616 131316 158672
rect 131252 158612 131316 158616
rect 132356 158672 132420 158676
rect 132356 158616 132406 158672
rect 132406 158616 132420 158672
rect 132356 158612 132420 158616
rect 133460 158672 133524 158676
rect 133460 158616 133510 158672
rect 133510 158616 133524 158672
rect 133460 158612 133524 158616
rect 138612 158612 138676 158676
rect 159220 158612 159284 158676
rect 168236 158672 168300 158676
rect 168236 158616 168286 158672
rect 168286 158616 168300 158672
rect 168236 158612 168300 158616
rect 188660 158672 188724 158676
rect 188660 158616 188710 158672
rect 188710 158616 188724 158672
rect 188660 158612 188724 158616
rect 205956 158672 206020 158676
rect 205956 158616 206006 158672
rect 206006 158616 206020 158672
rect 205956 158612 206020 158616
rect 315804 158612 315868 158676
rect 317092 158672 317156 158676
rect 317092 158616 317106 158672
rect 317106 158616 317156 158672
rect 317092 158612 317156 158616
rect 319484 158672 319548 158676
rect 319484 158616 319498 158672
rect 319498 158616 319548 158672
rect 319484 158612 319548 158616
rect 320588 158672 320652 158676
rect 320588 158616 320602 158672
rect 320602 158616 320652 158672
rect 320588 158612 320652 158616
rect 321692 158672 321756 158676
rect 321692 158616 321706 158672
rect 321706 158616 321756 158672
rect 321692 158612 321756 158616
rect 323164 158672 323228 158676
rect 323164 158616 323178 158672
rect 323178 158616 323228 158672
rect 323164 158612 323228 158616
rect 327580 158672 327644 158676
rect 327580 158616 327594 158672
rect 327594 158616 327644 158672
rect 327580 158612 327644 158616
rect 328316 158672 328380 158676
rect 328316 158616 328330 158672
rect 328330 158616 328380 158672
rect 328316 158612 328380 158616
rect 329972 158672 330036 158676
rect 329972 158616 329986 158672
rect 329986 158616 330036 158672
rect 329972 158612 330036 158616
rect 330708 158612 330772 158676
rect 331260 158672 331324 158676
rect 331260 158616 331274 158672
rect 331274 158616 331324 158672
rect 331260 158612 331324 158616
rect 332364 158672 332428 158676
rect 332364 158616 332378 158672
rect 332378 158616 332428 158672
rect 332364 158612 332428 158616
rect 333652 158672 333716 158676
rect 333652 158616 333666 158672
rect 333666 158616 333716 158672
rect 333652 158612 333716 158616
rect 334572 158672 334636 158676
rect 334572 158616 334586 158672
rect 334586 158616 334636 158672
rect 334572 158612 334636 158616
rect 335860 158672 335924 158676
rect 335860 158616 335874 158672
rect 335874 158616 335924 158672
rect 335860 158612 335924 158616
rect 336044 158672 336108 158676
rect 336044 158616 336058 158672
rect 336058 158616 336108 158672
rect 336044 158612 336108 158616
rect 336964 158672 337028 158676
rect 336964 158616 336978 158672
rect 336978 158616 337028 158672
rect 336964 158612 337028 158616
rect 338436 158672 338500 158676
rect 338436 158616 338450 158672
rect 338450 158616 338500 158672
rect 338436 158612 338500 158616
rect 339356 158672 339420 158676
rect 339356 158616 339370 158672
rect 339370 158616 339420 158672
rect 339356 158612 339420 158616
rect 341012 158672 341076 158676
rect 341012 158616 341026 158672
rect 341026 158616 341076 158672
rect 341012 158612 341076 158616
rect 343588 158672 343652 158676
rect 343588 158616 343602 158672
rect 343602 158616 343652 158672
rect 343588 158612 343652 158616
rect 347636 158672 347700 158676
rect 347636 158616 347650 158672
rect 347650 158616 347700 158672
rect 347636 158612 347700 158616
rect 354444 158672 354508 158676
rect 354444 158616 354458 158672
rect 354458 158616 354508 158672
rect 354444 158612 354508 158616
rect 355732 158612 355796 158676
rect 357020 158672 357084 158676
rect 357020 158616 357034 158672
rect 357034 158616 357084 158672
rect 357020 158612 357084 158616
rect 363460 158672 363524 158676
rect 363460 158616 363474 158672
rect 363474 158616 363524 158672
rect 363460 158612 363524 158616
rect 371004 158672 371068 158676
rect 371004 158616 371018 158672
rect 371018 158616 371068 158672
rect 371004 158612 371068 158616
rect 373396 158672 373460 158676
rect 373396 158616 373446 158672
rect 373446 158616 373460 158672
rect 373396 158612 373460 158616
rect 375972 158672 376036 158676
rect 375972 158616 376022 158672
rect 376022 158616 376036 158672
rect 375972 158612 376036 158616
rect 378548 158672 378612 158676
rect 378548 158616 378598 158672
rect 378598 158616 378612 158672
rect 378548 158612 378612 158616
rect 380940 158672 381004 158676
rect 380940 158616 380990 158672
rect 380990 158616 381004 158672
rect 380940 158612 381004 158616
rect 383516 158672 383580 158676
rect 383516 158616 383566 158672
rect 383566 158616 383580 158672
rect 383516 158612 383580 158616
rect 385908 158672 385972 158676
rect 385908 158616 385958 158672
rect 385958 158616 385972 158672
rect 385908 158612 385972 158616
rect 388484 158672 388548 158676
rect 388484 158616 388534 158672
rect 388534 158616 388548 158672
rect 388484 158612 388548 158616
rect 391060 158612 391124 158676
rect 393452 158612 393516 158676
rect 395844 158672 395908 158676
rect 395844 158616 395894 158672
rect 395894 158616 395908 158672
rect 395844 158612 395908 158616
rect 398420 158672 398484 158676
rect 398420 158616 398470 158672
rect 398470 158616 398484 158672
rect 398420 158612 398484 158616
rect 400996 158672 401060 158676
rect 400996 158616 401046 158672
rect 401046 158616 401060 158672
rect 400996 158612 401060 158616
rect 403388 158612 403452 158676
rect 405964 158612 406028 158676
rect 135852 158536 135916 158540
rect 135852 158480 135902 158536
rect 135902 158480 135916 158536
rect 135852 158476 135916 158480
rect 136956 158536 137020 158540
rect 136956 158480 137006 158536
rect 137006 158480 137020 158536
rect 136956 158476 137020 158480
rect 138060 158476 138124 158540
rect 139532 158476 139596 158540
rect 158116 158476 158180 158540
rect 358124 158476 358188 158540
rect 183508 158340 183572 158404
rect 185900 158400 185964 158404
rect 185900 158344 185950 158400
rect 185950 158344 185964 158400
rect 185900 158340 185964 158344
rect 193444 158340 193508 158404
rect 123156 158204 123220 158268
rect 134564 158264 134628 158268
rect 134564 158208 134614 158264
rect 134614 158208 134628 158264
rect 134564 158204 134628 158208
rect 141188 158204 141252 158268
rect 141740 158264 141804 158268
rect 141740 158208 141790 158264
rect 141790 158208 141804 158264
rect 141740 158204 141804 158208
rect 145972 158264 146036 158268
rect 145972 158208 146022 158264
rect 146022 158208 146036 158264
rect 145972 158204 146036 158208
rect 146340 158264 146404 158268
rect 146340 158208 146390 158264
rect 146390 158208 146404 158264
rect 146340 158204 146404 158208
rect 150940 158264 151004 158268
rect 150940 158208 150990 158264
rect 150990 158208 151004 158264
rect 150940 158204 151004 158208
rect 191052 158204 191116 158268
rect 195836 158264 195900 158268
rect 195836 158208 195886 158264
rect 195886 158208 195900 158264
rect 195836 158204 195900 158208
rect 328684 158340 328748 158404
rect 333468 158204 333532 158268
rect 338068 158264 338132 158268
rect 338068 158208 338118 158264
rect 338118 158208 338132 158264
rect 338068 158204 338132 158208
rect 343956 158264 344020 158268
rect 343956 158208 343970 158264
rect 343970 158208 344020 158264
rect 343956 158204 344020 158208
rect 348740 158264 348804 158268
rect 348740 158208 348754 158264
rect 348754 158208 348804 158264
rect 348740 158204 348804 158208
rect 353340 158264 353404 158268
rect 353340 158208 353354 158264
rect 353354 158208 353404 158264
rect 353340 158204 353404 158208
rect 117084 158068 117148 158132
rect 147628 158068 147692 158132
rect 170996 158068 171060 158132
rect 326476 158068 326540 158132
rect 140636 157992 140700 157996
rect 140636 157936 140686 157992
rect 140686 157936 140700 157992
rect 140636 157932 140700 157936
rect 142844 157932 142908 157996
rect 143580 157932 143644 157996
rect 318196 157932 318260 157996
rect 341748 157932 341812 157996
rect 345244 157932 345308 157996
rect 346348 157992 346412 157996
rect 346348 157936 346398 157992
rect 346398 157936 346412 157992
rect 346348 157932 346412 157936
rect 130700 157796 130764 157860
rect 283788 157796 283852 157860
rect 324268 157856 324332 157860
rect 324268 157800 324282 157856
rect 324282 157800 324332 157856
rect 324268 157796 324332 157800
rect 340644 157796 340708 157860
rect 342852 157796 342916 157860
rect 145236 157720 145300 157724
rect 145236 157664 145286 157720
rect 145286 157664 145300 157720
rect 145236 157660 145300 157664
rect 148364 157720 148428 157724
rect 148364 157664 148414 157720
rect 148414 157664 148428 157720
rect 148364 157660 148428 157664
rect 148732 157720 148796 157724
rect 148732 157664 148782 157720
rect 148782 157664 148796 157720
rect 148732 157660 148796 157664
rect 178540 157660 178604 157724
rect 283604 157660 283668 157724
rect 124260 157524 124324 157588
rect 155724 157584 155788 157588
rect 155724 157528 155774 157584
rect 155774 157528 155788 157584
rect 155724 157524 155788 157528
rect 200988 157584 201052 157588
rect 200988 157528 201038 157584
rect 201038 157528 201052 157584
rect 200988 157524 201052 157528
rect 203380 157584 203444 157588
rect 203380 157528 203430 157584
rect 203430 157528 203444 157584
rect 203380 157524 203444 157528
rect 359228 157524 359292 157588
rect 125364 157448 125428 157452
rect 125364 157392 125414 157448
rect 125414 157392 125428 157448
rect 125364 157388 125428 157392
rect 133644 157448 133708 157452
rect 133644 157392 133694 157448
rect 133694 157392 133708 157448
rect 133644 157388 133708 157392
rect 136036 157448 136100 157452
rect 136036 157392 136086 157448
rect 136086 157392 136100 157448
rect 136036 157388 136100 157392
rect 143948 157448 144012 157452
rect 143948 157392 143998 157448
rect 143998 157392 144012 157448
rect 143948 157388 144012 157392
rect 149836 157448 149900 157452
rect 149836 157392 149886 157448
rect 149886 157392 149900 157448
rect 149836 157388 149900 157392
rect 151308 157448 151372 157452
rect 151308 157392 151358 157448
rect 151358 157392 151372 157448
rect 151308 157388 151372 157392
rect 152228 157388 152292 157452
rect 153332 157388 153396 157452
rect 154436 157448 154500 157452
rect 154436 157392 154486 157448
rect 154486 157392 154500 157448
rect 154436 157388 154500 157392
rect 157012 157448 157076 157452
rect 157012 157392 157062 157448
rect 157062 157392 157076 157448
rect 157012 157388 157076 157392
rect 180932 157388 180996 157452
rect 198412 157448 198476 157452
rect 198412 157392 198462 157448
rect 198462 157392 198476 157448
rect 198412 157388 198476 157392
rect 295012 157448 295076 157452
rect 295012 157392 295062 157448
rect 295062 157392 295076 157448
rect 295012 157388 295076 157392
rect 325372 157388 325436 157452
rect 345980 157388 346044 157452
rect 349844 157448 349908 157452
rect 349844 157392 349858 157448
rect 349858 157392 349908 157448
rect 349844 157388 349908 157392
rect 351132 157448 351196 157452
rect 351132 157392 351146 157448
rect 351146 157392 351196 157448
rect 351132 157388 351196 157392
rect 352236 157448 352300 157452
rect 352236 157392 352250 157448
rect 352250 157392 352300 157448
rect 352236 157388 352300 157392
rect 290596 156708 290660 156772
rect 290780 156632 290844 156636
rect 290780 156576 290794 156632
rect 290794 156576 290844 156632
rect 290780 156572 290844 156576
rect 289492 155892 289556 155956
rect 289124 155756 289188 155820
rect 275324 154396 275388 154460
rect 275140 154260 275204 154324
rect 288940 153036 289004 153100
rect 284892 152356 284956 152420
rect 277532 148276 277596 148340
rect 279004 147596 279068 147660
rect 277164 141340 277228 141404
rect 278820 128964 278884 129028
rect 298324 80684 298388 80748
rect 296484 18532 296548 18596
rect 287652 9556 287716 9620
rect 286548 9420 286612 9484
rect 286732 9284 286796 9348
rect 292252 9148 292316 9212
rect 288020 9012 288084 9076
rect 287836 8876 287900 8940
rect 293540 8740 293604 8804
rect 297404 6836 297468 6900
rect 298508 6700 298572 6764
rect 282500 6564 282564 6628
rect 282684 6428 282748 6492
rect 295932 6292 295996 6356
rect 292436 6156 292500 6220
rect 297588 6020 297652 6084
rect 297956 4932 298020 4996
rect 297772 4796 297836 4860
rect 296300 3980 296364 4044
rect 439452 3980 439516 4044
rect 286916 3844 286980 3908
rect 296116 3708 296180 3772
rect 295196 3572 295260 3636
rect 437796 3572 437860 3636
rect 293724 3436 293788 3500
rect 437428 3436 437492 3500
rect 439084 3496 439148 3500
rect 439084 3440 439134 3496
rect 439134 3440 439148 3496
rect 439084 3436 439148 3440
rect 288204 3300 288268 3364
rect 437612 3300 437676 3364
rect 285076 3164 285140 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 245308 101414 245898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 245308 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 245308 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 245308 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 245308 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 245308 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 245308 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 245308 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 245308 137414 245898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 245308 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 245308 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 245308 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 245308 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 245308 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 245308 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 245308 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 245308 173414 245898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 245308 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 245308 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 245308 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 245308 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 245308 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 245308 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 245308 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 245308 209414 245898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 565308 218414 578898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 565308 222914 583398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 565308 227414 587898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 565308 231914 592398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 565308 236414 596898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 565308 240914 565398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 565308 245414 569898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 565308 249914 574398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 565308 254414 578898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 565308 258914 583398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 565308 263414 587898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 565308 267914 592398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 565308 272414 596898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 565308 276914 565398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 565308 281414 569898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 565308 285914 574398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 565308 290414 578898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 565308 294914 583398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 565308 299414 587898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 565308 303914 592398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 565308 308414 596898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 565308 312914 565398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 565308 317414 569898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 565308 321914 574398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 565308 326414 578898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 565308 330914 583398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 565308 335414 587898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 565308 339914 592398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 565308 344414 596898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 565308 348914 565398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 565308 353414 569898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 565308 357914 574398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 220272 547954 220620 547986
rect 220272 547718 220328 547954
rect 220564 547718 220620 547954
rect 220272 547634 220620 547718
rect 220272 547398 220328 547634
rect 220564 547398 220620 547634
rect 220272 547366 220620 547398
rect 356000 547954 356348 547986
rect 356000 547718 356056 547954
rect 356292 547718 356348 547954
rect 356000 547634 356348 547718
rect 356000 547398 356056 547634
rect 356292 547398 356348 547634
rect 356000 547366 356348 547398
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 220272 511954 220620 511986
rect 220272 511718 220328 511954
rect 220564 511718 220620 511954
rect 220272 511634 220620 511718
rect 220272 511398 220328 511634
rect 220564 511398 220620 511634
rect 220272 511366 220620 511398
rect 356000 511954 356348 511986
rect 356000 511718 356056 511954
rect 356292 511718 356348 511954
rect 356000 511634 356348 511718
rect 356000 511398 356056 511634
rect 356292 511398 356348 511634
rect 356000 511366 356348 511398
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 236056 479770 236116 480080
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 235950 479710 236116 479770
rect 237054 479710 237204 479770
rect 238158 479710 238292 479770
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 241768 479710 241898 479770
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 245308 213914 250398
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 245308 218414 254898
rect 222294 475954 222914 478000
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 245308 222914 259398
rect 226794 444454 227414 478000
rect 235950 476373 236010 479710
rect 235947 476372 236013 476373
rect 235947 476308 235948 476372
rect 236012 476308 236013 476372
rect 235947 476307 236013 476308
rect 237054 476237 237114 479710
rect 238158 476237 238218 479710
rect 239630 476781 239690 479710
rect 239627 476780 239693 476781
rect 239627 476716 239628 476780
rect 239692 476716 239693 476780
rect 239627 476715 239693 476716
rect 240550 476237 240610 479710
rect 241838 476237 241898 479710
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244290 479770
rect 243126 476917 243186 479710
rect 243123 476916 243189 476917
rect 243123 476852 243124 476916
rect 243188 476852 243189 476916
rect 243123 476851 243189 476852
rect 244230 476373 244290 479710
rect 245334 479710 245500 479770
rect 246438 479710 246588 479770
rect 247542 479710 247676 479770
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 250064 479710 250178 479770
rect 245334 476509 245394 479710
rect 245331 476508 245397 476509
rect 245331 476444 245332 476508
rect 245396 476444 245397 476508
rect 245331 476443 245397 476444
rect 244227 476372 244293 476373
rect 244227 476308 244228 476372
rect 244292 476308 244293 476372
rect 244227 476307 244293 476308
rect 246438 476237 246498 479710
rect 247542 476237 247602 479710
rect 248278 476917 248338 479710
rect 248275 476916 248341 476917
rect 248275 476852 248276 476916
rect 248340 476852 248341 476916
rect 248275 476851 248341 476852
rect 248646 476373 248706 479710
rect 248643 476372 248709 476373
rect 248643 476308 248644 476372
rect 248708 476308 248709 476372
rect 248643 476307 248709 476308
rect 250118 476237 250178 479710
rect 250670 479710 250804 479770
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 251288 479710 251466 479770
rect 250670 477325 250730 479710
rect 250667 477324 250733 477325
rect 250667 477260 250668 477324
rect 250732 477260 250733 477324
rect 250667 477259 250733 477260
rect 251406 476237 251466 479710
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 252326 476373 252386 479710
rect 252323 476372 252389 476373
rect 252323 476308 252324 476372
rect 252388 476308 252389 476372
rect 252323 476307 252389 476308
rect 253430 476237 253490 479710
rect 253614 476917 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 258496 479770 258556 480080
rect 256048 479710 256250 479770
rect 257000 479710 257170 479770
rect 253611 476916 253677 476917
rect 253611 476852 253612 476916
rect 253676 476852 253677 476916
rect 253611 476851 253677 476852
rect 254534 476373 254594 479710
rect 254531 476372 254597 476373
rect 254531 476308 254532 476372
rect 254596 476308 254597 476372
rect 254531 476307 254597 476308
rect 255822 476237 255882 479710
rect 256190 476917 256250 479710
rect 256187 476916 256253 476917
rect 256187 476852 256188 476916
rect 256252 476852 256253 476916
rect 256187 476851 256253 476852
rect 257110 476781 257170 479710
rect 257846 479710 258148 479770
rect 258398 479710 258556 479770
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 259448 479710 259562 479770
rect 260672 479710 260850 479770
rect 257846 477050 257906 479710
rect 258027 477052 258093 477053
rect 258027 477050 258028 477052
rect 257846 476990 258028 477050
rect 258027 476988 258028 476990
rect 258092 476988 258093 477052
rect 258027 476987 258093 476988
rect 257107 476780 257173 476781
rect 257107 476716 257108 476780
rect 257172 476716 257173 476780
rect 257107 476715 257173 476716
rect 258398 476645 258458 479710
rect 258395 476644 258461 476645
rect 258395 476580 258396 476644
rect 258460 476580 258461 476644
rect 258395 476579 258461 476580
rect 259502 476237 259562 479710
rect 260790 476373 260850 479710
rect 260974 479710 261140 479770
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 263528 479710 263610 479770
rect 260974 476645 261034 479710
rect 260971 476644 261037 476645
rect 260971 476580 260972 476644
rect 261036 476580 261037 476644
rect 260971 476579 261037 476580
rect 260787 476372 260853 476373
rect 260787 476308 260788 476372
rect 260852 476308 260853 476372
rect 260787 476307 260853 476308
rect 261710 476237 261770 479710
rect 262814 476509 262874 479710
rect 263550 476781 263610 479710
rect 263918 479710 263996 479770
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 265296 479710 265450 479770
rect 263547 476780 263613 476781
rect 263547 476716 263548 476780
rect 263612 476716 263613 476780
rect 263547 476715 263613 476716
rect 262811 476508 262877 476509
rect 262811 476444 262812 476508
rect 262876 476444 262877 476508
rect 262811 476443 262877 476444
rect 263918 476373 263978 479710
rect 263915 476372 263981 476373
rect 263915 476308 263916 476372
rect 263980 476308 263981 476372
rect 263915 476307 263981 476308
rect 265390 476237 265450 479710
rect 265942 479710 266036 479770
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 266384 479710 266554 479770
rect 265942 476509 266002 479710
rect 265939 476508 266005 476509
rect 265939 476444 265940 476508
rect 266004 476444 266005 476508
rect 265939 476443 266005 476444
rect 266494 476237 266554 479710
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 267598 476373 267658 479710
rect 268334 477325 268394 479710
rect 268331 477324 268397 477325
rect 268331 477260 268332 477324
rect 268396 477260 268397 477324
rect 268331 477259 268397 477260
rect 267595 476372 267661 476373
rect 267595 476308 267596 476372
rect 267660 476308 267661 476372
rect 267595 476307 267661 476308
rect 268702 476237 268762 479710
rect 269806 476237 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 271144 479710 271338 479770
rect 270910 477053 270970 479710
rect 270907 477052 270973 477053
rect 270907 476988 270908 477052
rect 270972 476988 270973 477052
rect 270907 476987 270973 476988
rect 271278 476237 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273486 479710 273652 479770
rect 274406 479710 274468 479770
rect 275768 479770 275828 480080
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 275768 479710 275938 479770
rect 276040 479710 276122 479770
rect 272198 476237 272258 479710
rect 273302 476237 273362 479710
rect 273486 476373 273546 479710
rect 274406 476373 274466 479710
rect 273483 476372 273549 476373
rect 273483 476308 273484 476372
rect 273548 476308 273549 476372
rect 273483 476307 273549 476308
rect 274403 476372 274469 476373
rect 274403 476308 274404 476372
rect 274468 476308 274469 476372
rect 274403 476307 274469 476308
rect 275878 476237 275938 479710
rect 276062 476645 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276059 476644 276125 476645
rect 276059 476580 276060 476644
rect 276124 476580 276125 476644
rect 276059 476579 276125 476580
rect 276982 476237 277042 479710
rect 278086 476237 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 279168 479710 279250 479770
rect 278454 476917 278514 479710
rect 278451 476916 278517 476917
rect 278451 476852 278452 476916
rect 278516 476852 278517 476916
rect 278451 476851 278517 476852
rect 279190 476237 279250 479710
rect 280846 479710 280996 479770
rect 283422 479710 283580 479770
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 293448 479770 293508 480080
rect 285968 479710 286058 479770
rect 280846 476237 280906 479710
rect 283422 476237 283482 479710
rect 285998 476237 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293358 479710 293508 479770
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 288206 476237 288266 479710
rect 290966 476237 291026 479710
rect 293358 476237 293418 479710
rect 295934 476237 295994 479710
rect 298510 476237 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305870 479710 306020 479770
rect 308446 479710 308604 479770
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 318472 479770 318532 480080
rect 310992 479710 311082 479770
rect 300902 476237 300962 479710
rect 303478 476917 303538 479710
rect 305870 477053 305930 479710
rect 308446 477053 308506 479710
rect 305867 477052 305933 477053
rect 305867 476988 305868 477052
rect 305932 476988 305933 477052
rect 305867 476987 305933 476988
rect 308443 477052 308509 477053
rect 308443 476988 308444 477052
rect 308508 476988 308509 477052
rect 308443 476987 308509 476988
rect 311022 476917 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318382 479710 318532 479770
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 325952 479770 326012 480080
rect 320920 479710 321018 479770
rect 303475 476916 303541 476917
rect 303475 476852 303476 476916
rect 303540 476852 303541 476916
rect 303475 476851 303541 476852
rect 311019 476916 311085 476917
rect 311019 476852 311020 476916
rect 311084 476852 311085 476916
rect 311019 476851 311085 476852
rect 313414 476509 313474 479710
rect 315806 476509 315866 479710
rect 313411 476508 313477 476509
rect 313411 476444 313412 476508
rect 313476 476444 313477 476508
rect 313411 476443 313477 476444
rect 315803 476508 315869 476509
rect 315803 476444 315804 476508
rect 315868 476444 315869 476508
rect 315803 476443 315869 476444
rect 318382 476373 318442 479710
rect 320958 476373 321018 479710
rect 323350 479710 323428 479770
rect 325926 479710 326012 479770
rect 323350 476917 323410 479710
rect 325926 476917 325986 479710
rect 323347 476916 323413 476917
rect 323347 476852 323348 476916
rect 323412 476852 323413 476916
rect 323347 476851 323413 476852
rect 325923 476916 325989 476917
rect 325923 476852 325924 476916
rect 325988 476852 325989 476916
rect 325923 476851 325989 476852
rect 318379 476372 318445 476373
rect 318379 476308 318380 476372
rect 318444 476308 318445 476372
rect 318379 476307 318445 476308
rect 320955 476372 321021 476373
rect 320955 476308 320956 476372
rect 321020 476308 321021 476372
rect 320955 476307 321021 476308
rect 237051 476236 237117 476237
rect 237051 476172 237052 476236
rect 237116 476172 237117 476236
rect 237051 476171 237117 476172
rect 238155 476236 238221 476237
rect 238155 476172 238156 476236
rect 238220 476172 238221 476236
rect 238155 476171 238221 476172
rect 240547 476236 240613 476237
rect 240547 476172 240548 476236
rect 240612 476172 240613 476236
rect 240547 476171 240613 476172
rect 241835 476236 241901 476237
rect 241835 476172 241836 476236
rect 241900 476172 241901 476236
rect 241835 476171 241901 476172
rect 246435 476236 246501 476237
rect 246435 476172 246436 476236
rect 246500 476172 246501 476236
rect 246435 476171 246501 476172
rect 247539 476236 247605 476237
rect 247539 476172 247540 476236
rect 247604 476172 247605 476236
rect 247539 476171 247605 476172
rect 250115 476236 250181 476237
rect 250115 476172 250116 476236
rect 250180 476172 250181 476236
rect 250115 476171 250181 476172
rect 251403 476236 251469 476237
rect 251403 476172 251404 476236
rect 251468 476172 251469 476236
rect 251403 476171 251469 476172
rect 253427 476236 253493 476237
rect 253427 476172 253428 476236
rect 253492 476172 253493 476236
rect 253427 476171 253493 476172
rect 255819 476236 255885 476237
rect 255819 476172 255820 476236
rect 255884 476172 255885 476236
rect 255819 476171 255885 476172
rect 259499 476236 259565 476237
rect 259499 476172 259500 476236
rect 259564 476172 259565 476236
rect 259499 476171 259565 476172
rect 261707 476236 261773 476237
rect 261707 476172 261708 476236
rect 261772 476172 261773 476236
rect 261707 476171 261773 476172
rect 265387 476236 265453 476237
rect 265387 476172 265388 476236
rect 265452 476172 265453 476236
rect 265387 476171 265453 476172
rect 266491 476236 266557 476237
rect 266491 476172 266492 476236
rect 266556 476172 266557 476236
rect 266491 476171 266557 476172
rect 268699 476236 268765 476237
rect 268699 476172 268700 476236
rect 268764 476172 268765 476236
rect 268699 476171 268765 476172
rect 269803 476236 269869 476237
rect 269803 476172 269804 476236
rect 269868 476172 269869 476236
rect 269803 476171 269869 476172
rect 271275 476236 271341 476237
rect 271275 476172 271276 476236
rect 271340 476172 271341 476236
rect 271275 476171 271341 476172
rect 272195 476236 272261 476237
rect 272195 476172 272196 476236
rect 272260 476172 272261 476236
rect 272195 476171 272261 476172
rect 273299 476236 273365 476237
rect 273299 476172 273300 476236
rect 273364 476172 273365 476236
rect 273299 476171 273365 476172
rect 275875 476236 275941 476237
rect 275875 476172 275876 476236
rect 275940 476172 275941 476236
rect 275875 476171 275941 476172
rect 276979 476236 277045 476237
rect 276979 476172 276980 476236
rect 277044 476172 277045 476236
rect 276979 476171 277045 476172
rect 278083 476236 278149 476237
rect 278083 476172 278084 476236
rect 278148 476172 278149 476236
rect 278083 476171 278149 476172
rect 279187 476236 279253 476237
rect 279187 476172 279188 476236
rect 279252 476172 279253 476236
rect 279187 476171 279253 476172
rect 280843 476236 280909 476237
rect 280843 476172 280844 476236
rect 280908 476172 280909 476236
rect 280843 476171 280909 476172
rect 283419 476236 283485 476237
rect 283419 476172 283420 476236
rect 283484 476172 283485 476236
rect 283419 476171 283485 476172
rect 285995 476236 286061 476237
rect 285995 476172 285996 476236
rect 286060 476172 286061 476236
rect 285995 476171 286061 476172
rect 288203 476236 288269 476237
rect 288203 476172 288204 476236
rect 288268 476172 288269 476236
rect 288203 476171 288269 476172
rect 290963 476236 291029 476237
rect 290963 476172 290964 476236
rect 291028 476172 291029 476236
rect 290963 476171 291029 476172
rect 293355 476236 293421 476237
rect 293355 476172 293356 476236
rect 293420 476172 293421 476236
rect 293355 476171 293421 476172
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 298507 476236 298573 476237
rect 298507 476172 298508 476236
rect 298572 476172 298573 476236
rect 298507 476171 298573 476172
rect 300899 476236 300965 476237
rect 300899 476172 300900 476236
rect 300964 476172 300965 476236
rect 300899 476171 300965 476172
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 445608 362414 470898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 249568 439954 249888 439986
rect 249568 439718 249610 439954
rect 249846 439718 249888 439954
rect 249568 439634 249888 439718
rect 249568 439398 249610 439634
rect 249846 439398 249888 439634
rect 249568 439366 249888 439398
rect 280288 439954 280608 439986
rect 280288 439718 280330 439954
rect 280566 439718 280608 439954
rect 280288 439634 280608 439718
rect 280288 439398 280330 439634
rect 280566 439398 280608 439634
rect 280288 439366 280608 439398
rect 311008 439954 311328 439986
rect 311008 439718 311050 439954
rect 311286 439718 311328 439954
rect 311008 439634 311328 439718
rect 311008 439398 311050 439634
rect 311286 439398 311328 439634
rect 311008 439366 311328 439398
rect 341728 439954 342048 439986
rect 341728 439718 341770 439954
rect 342006 439718 342048 439954
rect 341728 439634 342048 439718
rect 341728 439398 341770 439634
rect 342006 439398 342048 439634
rect 341728 439366 342048 439398
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 234208 435454 234528 435486
rect 234208 435218 234250 435454
rect 234486 435218 234528 435454
rect 234208 435134 234528 435218
rect 234208 434898 234250 435134
rect 234486 434898 234528 435134
rect 234208 434866 234528 434898
rect 264928 435454 265248 435486
rect 264928 435218 264970 435454
rect 265206 435218 265248 435454
rect 264928 435134 265248 435218
rect 264928 434898 264970 435134
rect 265206 434898 265248 435134
rect 264928 434866 265248 434898
rect 295648 435454 295968 435486
rect 295648 435218 295690 435454
rect 295926 435218 295968 435454
rect 295648 435134 295968 435218
rect 295648 434898 295690 435134
rect 295926 434898 295968 435134
rect 295648 434866 295968 434898
rect 326368 435454 326688 435486
rect 326368 435218 326410 435454
rect 326646 435218 326688 435454
rect 326368 435134 326688 435218
rect 326368 434898 326410 435134
rect 326646 434898 326688 435134
rect 326368 434866 326688 434898
rect 357088 435454 357408 435486
rect 357088 435218 357130 435454
rect 357366 435218 357408 435454
rect 357088 435134 357408 435218
rect 357088 434898 357130 435134
rect 357366 434898 357408 435134
rect 357088 434866 357408 434898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 249568 403954 249888 403986
rect 249568 403718 249610 403954
rect 249846 403718 249888 403954
rect 249568 403634 249888 403718
rect 249568 403398 249610 403634
rect 249846 403398 249888 403634
rect 249568 403366 249888 403398
rect 280288 403954 280608 403986
rect 280288 403718 280330 403954
rect 280566 403718 280608 403954
rect 280288 403634 280608 403718
rect 280288 403398 280330 403634
rect 280566 403398 280608 403634
rect 280288 403366 280608 403398
rect 311008 403954 311328 403986
rect 311008 403718 311050 403954
rect 311286 403718 311328 403954
rect 311008 403634 311328 403718
rect 311008 403398 311050 403634
rect 311286 403398 311328 403634
rect 311008 403366 311328 403398
rect 341728 403954 342048 403986
rect 341728 403718 341770 403954
rect 342006 403718 342048 403954
rect 341728 403634 342048 403718
rect 341728 403398 341770 403634
rect 342006 403398 342048 403634
rect 341728 403366 342048 403398
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 234208 399454 234528 399486
rect 234208 399218 234250 399454
rect 234486 399218 234528 399454
rect 234208 399134 234528 399218
rect 234208 398898 234250 399134
rect 234486 398898 234528 399134
rect 234208 398866 234528 398898
rect 264928 399454 265248 399486
rect 264928 399218 264970 399454
rect 265206 399218 265248 399454
rect 264928 399134 265248 399218
rect 264928 398898 264970 399134
rect 265206 398898 265248 399134
rect 264928 398866 265248 398898
rect 295648 399454 295968 399486
rect 295648 399218 295690 399454
rect 295926 399218 295968 399454
rect 295648 399134 295968 399218
rect 295648 398898 295690 399134
rect 295926 398898 295968 399134
rect 295648 398866 295968 398898
rect 326368 399454 326688 399486
rect 326368 399218 326410 399454
rect 326646 399218 326688 399454
rect 326368 399134 326688 399218
rect 326368 398898 326410 399134
rect 326646 398898 326688 399134
rect 326368 398866 326688 398898
rect 357088 399454 357408 399486
rect 357088 399218 357130 399454
rect 357366 399218 357408 399454
rect 357088 399134 357408 399218
rect 357088 398898 357130 399134
rect 357366 398898 357408 399134
rect 357088 398866 357408 398898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 249568 367954 249888 367986
rect 249568 367718 249610 367954
rect 249846 367718 249888 367954
rect 249568 367634 249888 367718
rect 249568 367398 249610 367634
rect 249846 367398 249888 367634
rect 249568 367366 249888 367398
rect 280288 367954 280608 367986
rect 280288 367718 280330 367954
rect 280566 367718 280608 367954
rect 280288 367634 280608 367718
rect 280288 367398 280330 367634
rect 280566 367398 280608 367634
rect 280288 367366 280608 367398
rect 311008 367954 311328 367986
rect 311008 367718 311050 367954
rect 311286 367718 311328 367954
rect 311008 367634 311328 367718
rect 311008 367398 311050 367634
rect 311286 367398 311328 367634
rect 311008 367366 311328 367398
rect 341728 367954 342048 367986
rect 341728 367718 341770 367954
rect 342006 367718 342048 367954
rect 341728 367634 342048 367718
rect 341728 367398 341770 367634
rect 342006 367398 342048 367634
rect 341728 367366 342048 367398
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 234208 363454 234528 363486
rect 234208 363218 234250 363454
rect 234486 363218 234528 363454
rect 234208 363134 234528 363218
rect 234208 362898 234250 363134
rect 234486 362898 234528 363134
rect 234208 362866 234528 362898
rect 264928 363454 265248 363486
rect 264928 363218 264970 363454
rect 265206 363218 265248 363454
rect 264928 363134 265248 363218
rect 264928 362898 264970 363134
rect 265206 362898 265248 363134
rect 264928 362866 265248 362898
rect 295648 363454 295968 363486
rect 295648 363218 295690 363454
rect 295926 363218 295968 363454
rect 295648 363134 295968 363218
rect 295648 362898 295690 363134
rect 295926 362898 295968 363134
rect 295648 362866 295968 362898
rect 326368 363454 326688 363486
rect 326368 363218 326410 363454
rect 326646 363218 326688 363454
rect 326368 363134 326688 363218
rect 326368 362898 326410 363134
rect 326646 362898 326688 363134
rect 326368 362866 326688 362898
rect 357088 363454 357408 363486
rect 357088 363218 357130 363454
rect 357366 363218 357408 363454
rect 357088 363134 357408 363218
rect 357088 362898 357130 363134
rect 357366 362898 357408 363134
rect 357088 362866 357408 362898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 249568 331954 249888 331986
rect 249568 331718 249610 331954
rect 249846 331718 249888 331954
rect 249568 331634 249888 331718
rect 249568 331398 249610 331634
rect 249846 331398 249888 331634
rect 249568 331366 249888 331398
rect 280288 331954 280608 331986
rect 280288 331718 280330 331954
rect 280566 331718 280608 331954
rect 280288 331634 280608 331718
rect 280288 331398 280330 331634
rect 280566 331398 280608 331634
rect 280288 331366 280608 331398
rect 311008 331954 311328 331986
rect 311008 331718 311050 331954
rect 311286 331718 311328 331954
rect 311008 331634 311328 331718
rect 311008 331398 311050 331634
rect 311286 331398 311328 331634
rect 311008 331366 311328 331398
rect 341728 331954 342048 331986
rect 341728 331718 341770 331954
rect 342006 331718 342048 331954
rect 341728 331634 342048 331718
rect 341728 331398 341770 331634
rect 342006 331398 342048 331634
rect 341728 331366 342048 331398
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 234208 327454 234528 327486
rect 234208 327218 234250 327454
rect 234486 327218 234528 327454
rect 234208 327134 234528 327218
rect 234208 326898 234250 327134
rect 234486 326898 234528 327134
rect 234208 326866 234528 326898
rect 264928 327454 265248 327486
rect 264928 327218 264970 327454
rect 265206 327218 265248 327454
rect 264928 327134 265248 327218
rect 264928 326898 264970 327134
rect 265206 326898 265248 327134
rect 264928 326866 265248 326898
rect 295648 327454 295968 327486
rect 295648 327218 295690 327454
rect 295926 327218 295968 327454
rect 295648 327134 295968 327218
rect 295648 326898 295690 327134
rect 295926 326898 295968 327134
rect 295648 326866 295968 326898
rect 326368 327454 326688 327486
rect 326368 327218 326410 327454
rect 326646 327218 326688 327454
rect 326368 327134 326688 327218
rect 326368 326898 326410 327134
rect 326646 326898 326688 327134
rect 326368 326866 326688 326898
rect 357088 327454 357408 327486
rect 357088 327218 357130 327454
rect 357366 327218 357408 327454
rect 357088 327134 357408 327218
rect 357088 326898 357130 327134
rect 357366 326898 357408 327134
rect 357088 326866 357408 326898
rect 282683 309092 282749 309093
rect 282683 309028 282684 309092
rect 282748 309028 282749 309092
rect 282683 309027 282749 309028
rect 282131 308820 282197 308821
rect 282131 308756 282132 308820
rect 282196 308756 282197 308820
rect 282131 308755 282197 308756
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 245308 227414 263898
rect 231294 304954 231914 308400
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 245308 231914 268398
rect 240294 277954 240914 308400
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 100272 223954 100620 223986
rect 100272 223718 100328 223954
rect 100564 223718 100620 223954
rect 100272 223634 100620 223718
rect 100272 223398 100328 223634
rect 100564 223398 100620 223634
rect 100272 223366 100620 223398
rect 236000 223954 236348 223986
rect 236000 223718 236056 223954
rect 236292 223718 236348 223954
rect 236000 223634 236348 223718
rect 236000 223398 236056 223634
rect 236292 223398 236348 223634
rect 236000 223366 236348 223398
rect 100952 219454 101300 219486
rect 100952 219218 101008 219454
rect 101244 219218 101300 219454
rect 100952 219134 101300 219218
rect 100952 218898 101008 219134
rect 101244 218898 101300 219134
rect 100952 218866 101300 218898
rect 235320 219454 235668 219486
rect 235320 219218 235376 219454
rect 235612 219218 235668 219454
rect 235320 219134 235668 219218
rect 235320 218898 235376 219134
rect 235612 218898 235668 219134
rect 235320 218866 235668 218898
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 100272 187954 100620 187986
rect 100272 187718 100328 187954
rect 100564 187718 100620 187954
rect 100272 187634 100620 187718
rect 100272 187398 100328 187634
rect 100564 187398 100620 187634
rect 100272 187366 100620 187398
rect 236000 187954 236348 187986
rect 236000 187718 236056 187954
rect 236292 187718 236348 187954
rect 236000 187634 236348 187718
rect 236000 187398 236056 187634
rect 236292 187398 236348 187634
rect 236000 187366 236348 187398
rect 100952 183454 101300 183486
rect 100952 183218 101008 183454
rect 101244 183218 101300 183454
rect 100952 183134 101300 183218
rect 100952 182898 101008 183134
rect 101244 182898 101300 183134
rect 100952 182866 101300 182898
rect 235320 183454 235668 183486
rect 235320 183218 235376 183454
rect 235612 183218 235668 183454
rect 235320 183134 235668 183218
rect 235320 182898 235376 183134
rect 235612 182898 235668 183134
rect 235320 182866 235668 182898
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 116056 159490 116116 160106
rect 117144 159490 117204 160106
rect 118232 159490 118292 160106
rect 116056 159430 116226 159490
rect 116166 158677 116226 159430
rect 117086 159430 117204 159490
rect 118190 159430 118292 159490
rect 119592 159490 119652 160106
rect 120544 159490 120604 160106
rect 121768 159490 121828 160106
rect 123128 159490 123188 160106
rect 124216 159490 124276 160106
rect 125440 159490 125500 160106
rect 126528 159490 126588 160106
rect 127616 159490 127676 160106
rect 119592 159430 119722 159490
rect 120544 159430 120642 159490
rect 121768 159430 121930 159490
rect 123128 159430 123218 159490
rect 124216 159430 124322 159490
rect 116163 158676 116229 158677
rect 116163 158612 116164 158676
rect 116228 158612 116229 158676
rect 116163 158611 116229 158612
rect 117086 158133 117146 159430
rect 118190 158677 118250 159430
rect 119662 158677 119722 159430
rect 120582 158677 120642 159430
rect 121870 158677 121930 159430
rect 118187 158676 118253 158677
rect 118187 158612 118188 158676
rect 118252 158612 118253 158676
rect 118187 158611 118253 158612
rect 119659 158676 119725 158677
rect 119659 158612 119660 158676
rect 119724 158612 119725 158676
rect 119659 158611 119725 158612
rect 120579 158676 120645 158677
rect 120579 158612 120580 158676
rect 120644 158612 120645 158676
rect 120579 158611 120645 158612
rect 121867 158676 121933 158677
rect 121867 158612 121868 158676
rect 121932 158612 121933 158676
rect 121867 158611 121933 158612
rect 123158 158269 123218 159430
rect 123155 158268 123221 158269
rect 123155 158204 123156 158268
rect 123220 158204 123221 158268
rect 123155 158203 123221 158204
rect 117083 158132 117149 158133
rect 117083 158068 117084 158132
rect 117148 158068 117149 158132
rect 117083 158067 117149 158068
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 138454 101414 158000
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 142954 105914 158000
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 147454 110414 158000
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 151954 114914 158000
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 156454 119414 158000
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 124954 123914 158000
rect 124262 157589 124322 159430
rect 125366 159430 125500 159490
rect 126470 159430 126588 159490
rect 127574 159430 127676 159490
rect 128296 159490 128356 160106
rect 128704 159490 128764 160106
rect 128296 159430 128370 159490
rect 124259 157588 124325 157589
rect 124259 157524 124260 157588
rect 124324 157524 124325 157588
rect 124259 157523 124325 157524
rect 125366 157453 125426 159430
rect 126470 158677 126530 159430
rect 127574 158677 127634 159430
rect 128310 159221 128370 159430
rect 128678 159430 128764 159490
rect 130064 159490 130124 160106
rect 130744 159490 130804 160106
rect 131288 159490 131348 160106
rect 132376 159490 132436 160106
rect 133464 159490 133524 160106
rect 130064 159430 130210 159490
rect 128307 159220 128373 159221
rect 128307 159156 128308 159220
rect 128372 159156 128373 159220
rect 128307 159155 128373 159156
rect 128678 158677 128738 159430
rect 130150 158677 130210 159430
rect 130702 159430 130804 159490
rect 131254 159430 131348 159490
rect 132358 159430 132436 159490
rect 133462 159430 133524 159490
rect 133600 159490 133660 160106
rect 134552 159490 134612 160106
rect 135912 159490 135972 160106
rect 136048 159490 136108 160106
rect 137000 159490 137060 160106
rect 138088 159490 138148 160106
rect 133600 159430 133706 159490
rect 134552 159430 134626 159490
rect 126467 158676 126533 158677
rect 126467 158612 126468 158676
rect 126532 158612 126533 158676
rect 126467 158611 126533 158612
rect 127571 158676 127637 158677
rect 127571 158612 127572 158676
rect 127636 158612 127637 158676
rect 127571 158611 127637 158612
rect 128675 158676 128741 158677
rect 128675 158612 128676 158676
rect 128740 158612 128741 158676
rect 128675 158611 128741 158612
rect 130147 158676 130213 158677
rect 130147 158612 130148 158676
rect 130212 158612 130213 158676
rect 130147 158611 130213 158612
rect 125363 157452 125429 157453
rect 125363 157388 125364 157452
rect 125428 157388 125429 157452
rect 125363 157387 125429 157388
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 129454 128414 158000
rect 130702 157861 130762 159430
rect 131254 158677 131314 159430
rect 132358 158677 132418 159430
rect 133462 158677 133522 159430
rect 131251 158676 131317 158677
rect 131251 158612 131252 158676
rect 131316 158612 131317 158676
rect 131251 158611 131317 158612
rect 132355 158676 132421 158677
rect 132355 158612 132356 158676
rect 132420 158612 132421 158676
rect 132355 158611 132421 158612
rect 133459 158676 133525 158677
rect 133459 158612 133460 158676
rect 133524 158612 133525 158676
rect 133459 158611 133525 158612
rect 130699 157860 130765 157861
rect 130699 157796 130700 157860
rect 130764 157796 130765 157860
rect 130699 157795 130765 157796
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 133954 132914 158000
rect 133646 157453 133706 159430
rect 134566 158269 134626 159430
rect 135854 159430 135972 159490
rect 136038 159430 136108 159490
rect 136958 159430 137060 159490
rect 138062 159430 138148 159490
rect 138496 159490 138556 160106
rect 139448 159490 139508 160106
rect 140672 159490 140732 160106
rect 138496 159430 138674 159490
rect 139448 159430 139594 159490
rect 135854 158541 135914 159430
rect 135851 158540 135917 158541
rect 135851 158476 135852 158540
rect 135916 158476 135917 158540
rect 135851 158475 135917 158476
rect 134563 158268 134629 158269
rect 134563 158204 134564 158268
rect 134628 158204 134629 158268
rect 134563 158203 134629 158204
rect 136038 157453 136098 159430
rect 136958 158541 137018 159430
rect 138062 158541 138122 159430
rect 138614 158677 138674 159430
rect 138611 158676 138677 158677
rect 138611 158612 138612 158676
rect 138676 158612 138677 158676
rect 138611 158611 138677 158612
rect 139534 158541 139594 159430
rect 140638 159430 140732 159490
rect 141080 159490 141140 160106
rect 141760 159490 141820 160106
rect 142848 159490 142908 160106
rect 141080 159430 141250 159490
rect 136955 158540 137021 158541
rect 136955 158476 136956 158540
rect 137020 158476 137021 158540
rect 136955 158475 137021 158476
rect 138059 158540 138125 158541
rect 138059 158476 138060 158540
rect 138124 158476 138125 158540
rect 138059 158475 138125 158476
rect 139531 158540 139597 158541
rect 139531 158476 139532 158540
rect 139596 158476 139597 158540
rect 139531 158475 139597 158476
rect 133643 157452 133709 157453
rect 133643 157388 133644 157452
rect 133708 157388 133709 157452
rect 133643 157387 133709 157388
rect 136035 157452 136101 157453
rect 136035 157388 136036 157452
rect 136100 157388 136101 157452
rect 136035 157387 136101 157388
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 138454 137414 158000
rect 140638 157997 140698 159430
rect 141190 158269 141250 159430
rect 141742 159430 141820 159490
rect 142846 159430 142908 159490
rect 143528 159490 143588 160106
rect 143936 159490 143996 160106
rect 145296 159490 145356 160106
rect 145976 159490 146036 160106
rect 146384 159490 146444 160106
rect 143528 159430 143642 159490
rect 143936 159430 144010 159490
rect 141742 158269 141802 159430
rect 141187 158268 141253 158269
rect 141187 158204 141188 158268
rect 141252 158204 141253 158268
rect 141187 158203 141253 158204
rect 141739 158268 141805 158269
rect 141739 158204 141740 158268
rect 141804 158204 141805 158268
rect 141739 158203 141805 158204
rect 140635 157996 140701 157997
rect 140635 157932 140636 157996
rect 140700 157932 140701 157996
rect 140635 157931 140701 157932
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 142954 141914 158000
rect 142846 157997 142906 159430
rect 143582 157997 143642 159430
rect 142843 157996 142909 157997
rect 142843 157932 142844 157996
rect 142908 157932 142909 157996
rect 142843 157931 142909 157932
rect 143579 157996 143645 157997
rect 143579 157932 143580 157996
rect 143644 157932 143645 157996
rect 143579 157931 143645 157932
rect 143950 157453 144010 159430
rect 145238 159430 145356 159490
rect 145974 159430 146036 159490
rect 146342 159430 146444 159490
rect 147608 159490 147668 160106
rect 148288 159490 148348 160106
rect 148696 159490 148756 160106
rect 149784 159490 149844 160106
rect 151008 159490 151068 160106
rect 147608 159430 147690 159490
rect 148288 159430 148426 159490
rect 148696 159430 148794 159490
rect 149784 159430 149898 159490
rect 145238 157725 145298 159430
rect 145974 158269 146034 159430
rect 146342 158269 146402 159430
rect 145971 158268 146037 158269
rect 145971 158204 145972 158268
rect 146036 158204 146037 158268
rect 145971 158203 146037 158204
rect 146339 158268 146405 158269
rect 146339 158204 146340 158268
rect 146404 158204 146405 158268
rect 146339 158203 146405 158204
rect 147630 158133 147690 159430
rect 147627 158132 147693 158133
rect 147627 158068 147628 158132
rect 147692 158068 147693 158132
rect 147627 158067 147693 158068
rect 145235 157724 145301 157725
rect 145235 157660 145236 157724
rect 145300 157660 145301 157724
rect 145235 157659 145301 157660
rect 143947 157452 144013 157453
rect 143947 157388 143948 157452
rect 144012 157388 144013 157452
rect 143947 157387 144013 157388
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 147454 146414 158000
rect 148366 157725 148426 159430
rect 148734 157725 148794 159430
rect 148363 157724 148429 157725
rect 148363 157660 148364 157724
rect 148428 157660 148429 157724
rect 148363 157659 148429 157660
rect 148731 157724 148797 157725
rect 148731 157660 148732 157724
rect 148796 157660 148797 157724
rect 148731 157659 148797 157660
rect 149838 157453 149898 159430
rect 150942 159430 151068 159490
rect 151144 159490 151204 160106
rect 152232 159490 152292 160106
rect 151144 159430 151370 159490
rect 150942 158269 151002 159430
rect 150939 158268 151005 158269
rect 150939 158204 150940 158268
rect 151004 158204 151005 158268
rect 150939 158203 151005 158204
rect 149835 157452 149901 157453
rect 149835 157388 149836 157452
rect 149900 157388 149901 157452
rect 149835 157387 149901 157388
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 151954 150914 158000
rect 151310 157453 151370 159430
rect 152230 159430 152292 159490
rect 153320 159490 153380 160106
rect 153592 159901 153652 160106
rect 153589 159900 153655 159901
rect 153589 159836 153590 159900
rect 153654 159836 153655 159900
rect 153589 159835 153655 159836
rect 154408 159490 154468 160106
rect 155768 159490 155828 160106
rect 156040 159901 156100 160106
rect 156037 159900 156103 159901
rect 156037 159836 156038 159900
rect 156102 159836 156103 159900
rect 156037 159835 156103 159836
rect 153320 159430 153394 159490
rect 154408 159430 154498 159490
rect 152230 157453 152290 159430
rect 153334 157453 153394 159430
rect 154438 157453 154498 159430
rect 155726 159430 155828 159490
rect 156992 159490 157052 160106
rect 158080 159490 158140 160106
rect 158488 159490 158548 160106
rect 156992 159430 157074 159490
rect 158080 159430 158178 159490
rect 151307 157452 151373 157453
rect 151307 157388 151308 157452
rect 151372 157388 151373 157452
rect 151307 157387 151373 157388
rect 152227 157452 152293 157453
rect 152227 157388 152228 157452
rect 152292 157388 152293 157452
rect 152227 157387 152293 157388
rect 153331 157452 153397 157453
rect 153331 157388 153332 157452
rect 153396 157388 153397 157452
rect 153331 157387 153397 157388
rect 154435 157452 154501 157453
rect 154435 157388 154436 157452
rect 154500 157388 154501 157452
rect 154435 157387 154501 157388
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 156454 155414 158000
rect 155726 157589 155786 159430
rect 155723 157588 155789 157589
rect 155723 157524 155724 157588
rect 155788 157524 155789 157588
rect 155723 157523 155789 157524
rect 157014 157453 157074 159430
rect 158118 158541 158178 159430
rect 158486 159430 158548 159490
rect 159168 159490 159228 160106
rect 160936 159901 160996 160106
rect 160933 159900 160999 159901
rect 160933 159836 160934 159900
rect 160998 159836 160999 159900
rect 160933 159835 160999 159836
rect 163520 159490 163580 160106
rect 165968 159629 166028 160106
rect 165965 159628 166031 159629
rect 165965 159564 165966 159628
rect 166030 159564 166031 159628
rect 165965 159563 166031 159564
rect 168280 159490 168340 160106
rect 171000 159490 171060 160106
rect 173448 159490 173508 160106
rect 175896 159901 175956 160106
rect 175893 159900 175959 159901
rect 175893 159836 175894 159900
rect 175958 159836 175959 159900
rect 175893 159835 175959 159836
rect 159168 159430 159282 159490
rect 163520 159430 163698 159490
rect 158486 158813 158546 159430
rect 158483 158812 158549 158813
rect 158483 158748 158484 158812
rect 158548 158748 158549 158812
rect 158483 158747 158549 158748
rect 159222 158677 159282 159430
rect 163638 158949 163698 159430
rect 168238 159430 168340 159490
rect 170998 159430 171060 159490
rect 173390 159430 173508 159490
rect 178480 159490 178540 160106
rect 180928 159490 180988 160106
rect 183512 159490 183572 160106
rect 185960 159490 186020 160106
rect 178480 159430 178602 159490
rect 180928 159430 180994 159490
rect 163635 158948 163701 158949
rect 163635 158884 163636 158948
rect 163700 158884 163701 158948
rect 163635 158883 163701 158884
rect 168238 158677 168298 159430
rect 159219 158676 159285 158677
rect 159219 158612 159220 158676
rect 159284 158612 159285 158676
rect 159219 158611 159285 158612
rect 168235 158676 168301 158677
rect 168235 158612 168236 158676
rect 168300 158612 168301 158676
rect 168235 158611 168301 158612
rect 158115 158540 158181 158541
rect 158115 158476 158116 158540
rect 158180 158476 158181 158540
rect 158115 158475 158181 158476
rect 170998 158133 171058 159430
rect 173390 159085 173450 159430
rect 173387 159084 173453 159085
rect 173387 159020 173388 159084
rect 173452 159020 173453 159084
rect 173387 159019 173453 159020
rect 170995 158132 171061 158133
rect 170995 158068 170996 158132
rect 171060 158068 171061 158132
rect 170995 158067 171061 158068
rect 157011 157452 157077 157453
rect 157011 157388 157012 157452
rect 157076 157388 157077 157452
rect 157011 157387 157077 157388
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 124954 159914 158000
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 129454 164414 158000
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 133954 168914 158000
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 138454 173414 158000
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 142954 177914 158000
rect 178542 157725 178602 159430
rect 178539 157724 178605 157725
rect 178539 157660 178540 157724
rect 178604 157660 178605 157724
rect 178539 157659 178605 157660
rect 180934 157453 180994 159430
rect 183510 159430 183572 159490
rect 185902 159430 186020 159490
rect 188544 159490 188604 160106
rect 190992 159490 191052 160106
rect 193440 159490 193500 160106
rect 195888 159490 195948 160106
rect 198472 159490 198532 160106
rect 188544 159430 188722 159490
rect 190992 159430 191114 159490
rect 193440 159430 193506 159490
rect 183510 158405 183570 159430
rect 185902 158405 185962 159430
rect 188662 158677 188722 159430
rect 188659 158676 188725 158677
rect 188659 158612 188660 158676
rect 188724 158612 188725 158676
rect 188659 158611 188725 158612
rect 183507 158404 183573 158405
rect 183507 158340 183508 158404
rect 183572 158340 183573 158404
rect 183507 158339 183573 158340
rect 185899 158404 185965 158405
rect 185899 158340 185900 158404
rect 185964 158340 185965 158404
rect 185899 158339 185965 158340
rect 191054 158269 191114 159430
rect 193446 158405 193506 159430
rect 195838 159430 195948 159490
rect 198414 159430 198532 159490
rect 200920 159490 200980 160106
rect 203368 159490 203428 160106
rect 205952 159490 206012 160106
rect 200920 159430 201050 159490
rect 203368 159430 203442 159490
rect 205952 159430 206018 159490
rect 193443 158404 193509 158405
rect 193443 158340 193444 158404
rect 193508 158340 193509 158404
rect 193443 158339 193509 158340
rect 195838 158269 195898 159430
rect 191051 158268 191117 158269
rect 191051 158204 191052 158268
rect 191116 158204 191117 158268
rect 191051 158203 191117 158204
rect 195835 158268 195901 158269
rect 195835 158204 195836 158268
rect 195900 158204 195901 158268
rect 195835 158203 195901 158204
rect 180931 157452 180997 157453
rect 180931 157388 180932 157452
rect 180996 157388 180997 157452
rect 180931 157387 180997 157388
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 147454 182414 158000
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 151954 186914 158000
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 156454 191414 158000
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 124954 195914 158000
rect 198414 157453 198474 159430
rect 198411 157452 198477 157453
rect 198411 157388 198412 157452
rect 198476 157388 198477 157452
rect 198411 157387 198477 157388
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 129454 200414 158000
rect 200990 157589 201050 159430
rect 203382 157589 203442 159430
rect 205958 158677 206018 159430
rect 205955 158676 206021 158677
rect 205955 158612 205956 158676
rect 206020 158612 206021 158676
rect 205955 158611 206021 158612
rect 200987 157588 201053 157589
rect 200987 157524 200988 157588
rect 201052 157524 201053 157588
rect 200987 157523 201053 157524
rect 203379 157588 203445 157589
rect 203379 157524 203380 157588
rect 203444 157524 203445 157588
rect 203379 157523 203445 157524
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 133954 204914 158000
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 138454 209414 158000
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 142954 213914 158000
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 151954 222914 158000
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 156454 227414 158000
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 124954 231914 158000
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 129454 236414 158000
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 282454 245414 308400
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 286954 249914 308400
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 291454 254414 308400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 295954 258914 308400
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 300454 263414 308400
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 304954 267914 308400
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 273454 272414 308400
rect 275323 303380 275389 303381
rect 275323 303316 275324 303380
rect 275388 303316 275389 303380
rect 275323 303315 275389 303316
rect 275139 303244 275205 303245
rect 275139 303180 275140 303244
rect 275204 303180 275205 303244
rect 275139 303179 275205 303180
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 275142 154325 275202 303179
rect 275326 154461 275386 303315
rect 276294 277954 276914 308400
rect 277347 308004 277413 308005
rect 277347 307940 277348 308004
rect 277412 307940 277413 308004
rect 277347 307939 277413 307940
rect 277350 302250 277410 307939
rect 277531 307868 277597 307869
rect 277531 307804 277532 307868
rect 277596 307804 277597 307868
rect 277531 307803 277597 307804
rect 278819 307868 278885 307869
rect 278819 307804 278820 307868
rect 278884 307804 278885 307868
rect 278819 307803 278885 307804
rect 279003 307868 279069 307869
rect 279003 307804 279004 307868
rect 279068 307804 279069 307868
rect 279003 307803 279069 307804
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 275323 154460 275389 154461
rect 275323 154396 275324 154460
rect 275388 154396 275389 154460
rect 275323 154395 275389 154396
rect 275139 154324 275205 154325
rect 275139 154260 275140 154324
rect 275204 154260 275205 154324
rect 275139 154259 275205 154260
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 133954 276914 169398
rect 277166 302190 277410 302250
rect 277166 141405 277226 302190
rect 277534 148341 277594 307803
rect 277531 148340 277597 148341
rect 277531 148276 277532 148340
rect 277596 148276 277597 148340
rect 277531 148275 277597 148276
rect 277163 141404 277229 141405
rect 277163 141340 277164 141404
rect 277228 141340 277229 141404
rect 277163 141339 277229 141340
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 278822 129029 278882 307803
rect 279006 147661 279066 307803
rect 280794 282454 281414 308400
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 279003 147660 279069 147661
rect 279003 147596 279004 147660
rect 279068 147596 279069 147660
rect 279003 147595 279069 147596
rect 280794 138454 281414 173898
rect 282134 158949 282194 308755
rect 282499 244900 282565 244901
rect 282499 244836 282500 244900
rect 282564 244836 282565 244900
rect 282499 244835 282565 244836
rect 282131 158948 282197 158949
rect 282131 158884 282132 158948
rect 282196 158884 282197 158948
rect 282131 158883 282197 158884
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 278819 129028 278885 129029
rect 278819 128964 278820 129028
rect 278884 128964 278885 129028
rect 278819 128963 278885 128964
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 282502 6629 282562 244835
rect 282499 6628 282565 6629
rect 282499 6564 282500 6628
rect 282564 6564 282565 6628
rect 282499 6563 282565 6564
rect 282686 6493 282746 309027
rect 283419 308956 283485 308957
rect 283419 308892 283420 308956
rect 283484 308892 283485 308956
rect 283419 308891 283485 308892
rect 283422 158813 283482 308891
rect 284707 308548 284773 308549
rect 284707 308484 284708 308548
rect 284772 308484 284773 308548
rect 284707 308483 284773 308484
rect 283787 306236 283853 306237
rect 283787 306172 283788 306236
rect 283852 306172 283853 306236
rect 283787 306171 283853 306172
rect 283603 306100 283669 306101
rect 283603 306036 283604 306100
rect 283668 306036 283669 306100
rect 283603 306035 283669 306036
rect 283419 158812 283485 158813
rect 283419 158748 283420 158812
rect 283484 158748 283485 158812
rect 283419 158747 283485 158748
rect 283606 157725 283666 306035
rect 283790 157861 283850 306171
rect 284710 159085 284770 308483
rect 284891 307868 284957 307869
rect 284891 307804 284892 307868
rect 284956 307804 284957 307868
rect 284891 307803 284957 307804
rect 284707 159084 284773 159085
rect 284707 159020 284708 159084
rect 284772 159020 284773 159084
rect 284707 159019 284773 159020
rect 283787 157860 283853 157861
rect 283787 157796 283788 157860
rect 283852 157796 283853 157860
rect 283787 157795 283853 157796
rect 283603 157724 283669 157725
rect 283603 157660 283604 157724
rect 283668 157660 283669 157724
rect 283603 157659 283669 157660
rect 284894 152421 284954 307803
rect 285294 286954 285914 308400
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285075 246260 285141 246261
rect 285075 246196 285076 246260
rect 285140 246196 285141 246260
rect 285075 246195 285141 246196
rect 284891 152420 284957 152421
rect 284891 152356 284892 152420
rect 284956 152356 284957 152420
rect 284891 152355 284957 152356
rect 282683 6492 282749 6493
rect 282683 6428 282684 6492
rect 282748 6428 282749 6492
rect 282683 6427 282749 6428
rect 285078 3229 285138 246195
rect 285294 214954 285914 250398
rect 289794 291454 290414 308400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 287651 248164 287717 248165
rect 287651 248100 287652 248164
rect 287716 248100 287717 248164
rect 287651 248099 287717 248100
rect 286915 248028 286981 248029
rect 286915 247964 286916 248028
rect 286980 247964 286981 248028
rect 286915 247963 286981 247964
rect 286547 247620 286613 247621
rect 286547 247556 286548 247620
rect 286612 247556 286613 247620
rect 286547 247555 286613 247556
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285075 3228 285141 3229
rect 285075 3164 285076 3228
rect 285140 3164 285141 3228
rect 285075 3163 285141 3164
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 -7066 285914 34398
rect 286550 9485 286610 247555
rect 286731 247076 286797 247077
rect 286731 247012 286732 247076
rect 286796 247012 286797 247076
rect 286731 247011 286797 247012
rect 286547 9484 286613 9485
rect 286547 9420 286548 9484
rect 286612 9420 286613 9484
rect 286547 9419 286613 9420
rect 286734 9349 286794 247011
rect 286731 9348 286797 9349
rect 286731 9284 286732 9348
rect 286796 9284 286797 9348
rect 286731 9283 286797 9284
rect 286918 3909 286978 247963
rect 287654 9621 287714 248099
rect 289491 247892 289557 247893
rect 289491 247828 289492 247892
rect 289556 247828 289557 247892
rect 289491 247827 289557 247828
rect 288203 247756 288269 247757
rect 288203 247692 288204 247756
rect 288268 247692 288269 247756
rect 288203 247691 288269 247692
rect 287835 247076 287901 247077
rect 287835 247012 287836 247076
rect 287900 247012 287901 247076
rect 287835 247011 287901 247012
rect 288019 247076 288085 247077
rect 288019 247012 288020 247076
rect 288084 247012 288085 247076
rect 288019 247011 288085 247012
rect 287651 9620 287717 9621
rect 287651 9556 287652 9620
rect 287716 9556 287717 9620
rect 287651 9555 287717 9556
rect 287838 8941 287898 247011
rect 288022 9077 288082 247011
rect 288019 9076 288085 9077
rect 288019 9012 288020 9076
rect 288084 9012 288085 9076
rect 288019 9011 288085 9012
rect 287835 8940 287901 8941
rect 287835 8876 287836 8940
rect 287900 8876 287901 8940
rect 287835 8875 287901 8876
rect 286915 3908 286981 3909
rect 286915 3844 286916 3908
rect 286980 3844 286981 3908
rect 286915 3843 286981 3844
rect 288206 3365 288266 247691
rect 288939 247076 289005 247077
rect 288939 247012 288940 247076
rect 289004 247012 289005 247076
rect 288939 247011 289005 247012
rect 289123 247076 289189 247077
rect 289123 247012 289124 247076
rect 289188 247012 289189 247076
rect 289123 247011 289189 247012
rect 288942 153101 289002 247011
rect 289126 155821 289186 247011
rect 289307 245036 289373 245037
rect 289307 244972 289308 245036
rect 289372 244972 289373 245036
rect 289307 244971 289373 244972
rect 289310 158813 289370 244971
rect 289307 158812 289373 158813
rect 289307 158748 289308 158812
rect 289372 158748 289373 158812
rect 289307 158747 289373 158748
rect 289494 155957 289554 247827
rect 289794 219454 290414 254898
rect 294294 295954 294914 308400
rect 297955 308276 298021 308277
rect 297955 308212 297956 308276
rect 298020 308212 298021 308276
rect 297955 308211 298021 308212
rect 297403 308140 297469 308141
rect 297403 308076 297404 308140
rect 297468 308076 297469 308140
rect 297403 308075 297469 308076
rect 296483 307868 296549 307869
rect 296483 307804 296484 307868
rect 296548 307804 296549 307868
rect 296483 307803 296549 307804
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 293539 247348 293605 247349
rect 293539 247284 293540 247348
rect 293604 247284 293605 247348
rect 293539 247283 293605 247284
rect 290595 247076 290661 247077
rect 290595 247012 290596 247076
rect 290660 247012 290661 247076
rect 290595 247011 290661 247012
rect 292251 247076 292317 247077
rect 292251 247012 292252 247076
rect 292316 247012 292317 247076
rect 292251 247011 292317 247012
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289491 155956 289557 155957
rect 289491 155892 289492 155956
rect 289556 155892 289557 155956
rect 289491 155891 289557 155892
rect 289123 155820 289189 155821
rect 289123 155756 289124 155820
rect 289188 155756 289189 155820
rect 289123 155755 289189 155756
rect 288939 153100 289005 153101
rect 288939 153036 288940 153100
rect 289004 153036 289005 153100
rect 288939 153035 289005 153036
rect 289794 147454 290414 182898
rect 290598 156773 290658 247011
rect 290779 245172 290845 245173
rect 290779 245108 290780 245172
rect 290844 245108 290845 245172
rect 290779 245107 290845 245108
rect 290595 156772 290661 156773
rect 290595 156708 290596 156772
rect 290660 156708 290661 156772
rect 290595 156707 290661 156708
rect 290782 156637 290842 245107
rect 291699 244356 291765 244357
rect 291699 244292 291700 244356
rect 291764 244292 291765 244356
rect 291699 244291 291765 244292
rect 291883 244356 291949 244357
rect 291883 244292 291884 244356
rect 291948 244292 291949 244356
rect 291883 244291 291949 244292
rect 291702 166293 291762 244291
rect 291886 196077 291946 244291
rect 291883 196076 291949 196077
rect 291883 196012 291884 196076
rect 291948 196012 291949 196076
rect 291883 196011 291949 196012
rect 291699 166292 291765 166293
rect 291699 166228 291700 166292
rect 291764 166228 291765 166292
rect 291699 166227 291765 166228
rect 290779 156636 290845 156637
rect 290779 156572 290780 156636
rect 290844 156572 290845 156636
rect 290779 156571 290845 156572
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 292254 9213 292314 247011
rect 292435 245308 292501 245309
rect 292435 245244 292436 245308
rect 292500 245244 292501 245308
rect 292435 245243 292501 245244
rect 292251 9212 292317 9213
rect 292251 9148 292252 9212
rect 292316 9148 292317 9212
rect 292251 9147 292317 9148
rect 292438 6221 292498 245243
rect 293171 244492 293237 244493
rect 293171 244428 293172 244492
rect 293236 244428 293237 244492
rect 293171 244427 293237 244428
rect 293174 158813 293234 244427
rect 293355 244356 293421 244357
rect 293355 244292 293356 244356
rect 293420 244292 293421 244356
rect 293355 244291 293421 244292
rect 293358 158949 293418 244291
rect 293355 158948 293421 158949
rect 293355 158884 293356 158948
rect 293420 158884 293421 158948
rect 293355 158883 293421 158884
rect 293171 158812 293237 158813
rect 293171 158748 293172 158812
rect 293236 158748 293237 158812
rect 293171 158747 293237 158748
rect 293542 8805 293602 247283
rect 293723 245172 293789 245173
rect 293723 245108 293724 245172
rect 293788 245108 293789 245172
rect 293723 245107 293789 245108
rect 293539 8804 293605 8805
rect 293539 8740 293540 8804
rect 293604 8740 293605 8804
rect 293539 8739 293605 8740
rect 292435 6220 292501 6221
rect 292435 6156 292436 6220
rect 292500 6156 292501 6220
rect 292435 6155 292501 6156
rect 293726 3501 293786 245107
rect 294294 223954 294914 259398
rect 295195 247484 295261 247485
rect 295195 247420 295196 247484
rect 295260 247420 295261 247484
rect 295195 247419 295261 247420
rect 295011 244764 295077 244765
rect 295011 244700 295012 244764
rect 295076 244700 295077 244764
rect 295011 244699 295077 244700
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 295014 157453 295074 244699
rect 295011 157452 295077 157453
rect 295011 157388 295012 157452
rect 295076 157388 295077 157452
rect 295011 157387 295077 157388
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 288203 3364 288269 3365
rect 288203 3300 288204 3364
rect 288268 3300 288269 3364
rect 288203 3299 288269 3300
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 293723 3500 293789 3501
rect 293723 3436 293724 3500
rect 293788 3436 293789 3500
rect 293723 3435 293789 3436
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 -1306 294914 7398
rect 295198 3637 295258 247419
rect 295931 245444 295997 245445
rect 295931 245380 295932 245444
rect 295996 245380 295997 245444
rect 295931 245379 295997 245380
rect 295934 6357 295994 245379
rect 296115 244764 296181 244765
rect 296115 244700 296116 244764
rect 296180 244700 296181 244764
rect 296115 244699 296181 244700
rect 295931 6356 295997 6357
rect 295931 6292 295932 6356
rect 295996 6292 295997 6356
rect 295931 6291 295997 6292
rect 296118 3773 296178 244699
rect 296299 244628 296365 244629
rect 296299 244564 296300 244628
rect 296364 244564 296365 244628
rect 296299 244563 296365 244564
rect 296302 4045 296362 244563
rect 296486 18597 296546 307803
rect 296483 18596 296549 18597
rect 296483 18532 296484 18596
rect 296548 18532 296549 18596
rect 296483 18531 296549 18532
rect 297406 6901 297466 308075
rect 297587 308004 297653 308005
rect 297587 307940 297588 308004
rect 297652 307940 297653 308004
rect 297587 307939 297653 307940
rect 297403 6900 297469 6901
rect 297403 6836 297404 6900
rect 297468 6836 297469 6900
rect 297403 6835 297469 6836
rect 297590 6085 297650 307939
rect 297771 307868 297837 307869
rect 297771 307804 297772 307868
rect 297836 307804 297837 307868
rect 297771 307803 297837 307804
rect 297587 6084 297653 6085
rect 297587 6020 297588 6084
rect 297652 6020 297653 6084
rect 297587 6019 297653 6020
rect 297774 4861 297834 307803
rect 297958 4997 298018 308211
rect 298323 308004 298389 308005
rect 298323 307940 298324 308004
rect 298388 307940 298389 308004
rect 298323 307939 298389 307940
rect 298139 244356 298205 244357
rect 298139 244292 298140 244356
rect 298204 244292 298205 244356
rect 298139 244291 298205 244292
rect 298142 187781 298202 244291
rect 298139 187780 298205 187781
rect 298139 187716 298140 187780
rect 298204 187716 298205 187780
rect 298139 187715 298205 187716
rect 298326 80749 298386 307939
rect 298507 307868 298573 307869
rect 298507 307804 298508 307868
rect 298572 307804 298573 307868
rect 298507 307803 298573 307804
rect 298323 80748 298389 80749
rect 298323 80684 298324 80748
rect 298388 80684 298389 80748
rect 298323 80683 298389 80684
rect 298510 6765 298570 307803
rect 298794 300454 299414 308400
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 245308 299414 263898
rect 303294 304954 303914 308400
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 245308 303914 268398
rect 316794 282454 317414 308400
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 245308 317414 245898
rect 321294 286954 321914 308400
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 245308 321914 250398
rect 325794 291454 326414 308400
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 245308 326414 254898
rect 330294 295954 330914 308400
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 245308 330914 259398
rect 334794 300454 335414 308400
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 245308 335414 263898
rect 339294 304954 339914 308400
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 245308 339914 268398
rect 352794 282454 353414 308400
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 245308 353414 245898
rect 357294 286954 357914 308400
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 245308 357914 250398
rect 361794 291454 362414 308400
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 245308 362414 254898
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 245308 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 245308 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 245308 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 245308 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 245308 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 245308 389414 245898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 245308 393914 250398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 245308 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 245308 402914 259398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 245308 407414 263898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 245308 411914 268398
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 245308 416414 272898
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 245308 420914 277398
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 245308 425414 245898
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 245308 429914 250398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 439451 302972 439517 302973
rect 439451 302908 439452 302972
rect 439516 302908 439517 302972
rect 439451 302907 439517 302908
rect 439083 298756 439149 298757
rect 439083 298692 439084 298756
rect 439148 298692 439149 298756
rect 439083 298691 439149 298692
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 437427 287740 437493 287741
rect 437427 287676 437428 287740
rect 437492 287676 437493 287740
rect 437427 287675 437493 287676
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 245308 434414 254898
rect 298691 244356 298757 244357
rect 298691 244292 298692 244356
rect 298756 244292 298757 244356
rect 298691 244291 298757 244292
rect 298694 158813 298754 244291
rect 300272 223954 300620 223986
rect 300272 223718 300328 223954
rect 300564 223718 300620 223954
rect 300272 223634 300620 223718
rect 300272 223398 300328 223634
rect 300564 223398 300620 223634
rect 300272 223366 300620 223398
rect 436000 223954 436348 223986
rect 436000 223718 436056 223954
rect 436292 223718 436348 223954
rect 436000 223634 436348 223718
rect 436000 223398 436056 223634
rect 436292 223398 436348 223634
rect 436000 223366 436348 223398
rect 300952 219454 301300 219486
rect 300952 219218 301008 219454
rect 301244 219218 301300 219454
rect 300952 219134 301300 219218
rect 300952 218898 301008 219134
rect 301244 218898 301300 219134
rect 300952 218866 301300 218898
rect 435320 219454 435668 219486
rect 435320 219218 435376 219454
rect 435612 219218 435668 219454
rect 435320 219134 435668 219218
rect 435320 218898 435376 219134
rect 435612 218898 435668 219134
rect 435320 218866 435668 218898
rect 300272 187954 300620 187986
rect 300272 187718 300328 187954
rect 300564 187718 300620 187954
rect 300272 187634 300620 187718
rect 300272 187398 300328 187634
rect 300564 187398 300620 187634
rect 300272 187366 300620 187398
rect 436000 187954 436348 187986
rect 436000 187718 436056 187954
rect 436292 187718 436348 187954
rect 436000 187634 436348 187718
rect 436000 187398 436056 187634
rect 436292 187398 436348 187634
rect 436000 187366 436348 187398
rect 300952 183454 301300 183486
rect 300952 183218 301008 183454
rect 301244 183218 301300 183454
rect 300952 183134 301300 183218
rect 300952 182898 301008 183134
rect 301244 182898 301300 183134
rect 300952 182866 301300 182898
rect 435320 183454 435668 183486
rect 435320 183218 435376 183454
rect 435612 183218 435668 183454
rect 435320 183134 435668 183218
rect 435320 182898 435376 183134
rect 435612 182898 435668 183134
rect 435320 182866 435668 182898
rect 316056 159490 316116 160106
rect 317144 159490 317204 160106
rect 318232 159490 318292 160106
rect 319592 159490 319652 160106
rect 315806 159430 316116 159490
rect 317094 159430 317204 159490
rect 318198 159430 318292 159490
rect 319486 159430 319652 159490
rect 320544 159490 320604 160106
rect 321768 159490 321828 160106
rect 320544 159430 320650 159490
rect 298691 158812 298757 158813
rect 298691 158748 298692 158812
rect 298756 158748 298757 158812
rect 298691 158747 298757 158748
rect 315806 158677 315866 159430
rect 317094 158677 317154 159430
rect 315803 158676 315869 158677
rect 315803 158612 315804 158676
rect 315868 158612 315869 158676
rect 315803 158611 315869 158612
rect 317091 158676 317157 158677
rect 317091 158612 317092 158676
rect 317156 158612 317157 158676
rect 317091 158611 317157 158612
rect 298794 156454 299414 158000
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298507 6764 298573 6765
rect 298507 6700 298508 6764
rect 298572 6700 298573 6764
rect 298507 6699 298573 6700
rect 297955 4996 298021 4997
rect 297955 4932 297956 4996
rect 298020 4932 298021 4996
rect 297955 4931 298021 4932
rect 297771 4860 297837 4861
rect 297771 4796 297772 4860
rect 297836 4796 297837 4860
rect 297771 4795 297837 4796
rect 296299 4044 296365 4045
rect 296299 3980 296300 4044
rect 296364 3980 296365 4044
rect 296299 3979 296365 3980
rect 296115 3772 296181 3773
rect 296115 3708 296116 3772
rect 296180 3708 296181 3772
rect 296115 3707 296181 3708
rect 295195 3636 295261 3637
rect 295195 3572 295196 3636
rect 295260 3572 295261 3636
rect 295195 3571 295261 3572
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 124954 303914 158000
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 129454 308414 158000
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 133954 312914 158000
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 138454 317414 158000
rect 318198 157997 318258 159430
rect 319486 158677 319546 159430
rect 320590 158677 320650 159430
rect 321694 159430 321828 159490
rect 323128 159490 323188 160106
rect 324216 159490 324276 160106
rect 325440 159490 325500 160106
rect 326528 159490 326588 160106
rect 327616 159490 327676 160106
rect 323128 159430 323226 159490
rect 324216 159430 324330 159490
rect 321694 158677 321754 159430
rect 323166 158677 323226 159430
rect 319483 158676 319549 158677
rect 319483 158612 319484 158676
rect 319548 158612 319549 158676
rect 319483 158611 319549 158612
rect 320587 158676 320653 158677
rect 320587 158612 320588 158676
rect 320652 158612 320653 158676
rect 320587 158611 320653 158612
rect 321691 158676 321757 158677
rect 321691 158612 321692 158676
rect 321756 158612 321757 158676
rect 321691 158611 321757 158612
rect 323163 158676 323229 158677
rect 323163 158612 323164 158676
rect 323228 158612 323229 158676
rect 323163 158611 323229 158612
rect 318195 157996 318261 157997
rect 318195 157932 318196 157996
rect 318260 157932 318261 157996
rect 318195 157931 318261 157932
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 142954 321914 158000
rect 324270 157861 324330 159430
rect 325374 159430 325500 159490
rect 326478 159430 326588 159490
rect 327582 159430 327676 159490
rect 328296 159490 328356 160106
rect 328704 159490 328764 160106
rect 330064 159490 330124 160106
rect 330744 159490 330804 160106
rect 331288 159490 331348 160106
rect 332376 159490 332436 160106
rect 328296 159430 328378 159490
rect 324267 157860 324333 157861
rect 324267 157796 324268 157860
rect 324332 157796 324333 157860
rect 324267 157795 324333 157796
rect 325374 157453 325434 159430
rect 326478 158133 326538 159430
rect 327582 158677 327642 159430
rect 328318 158677 328378 159430
rect 328686 159430 328764 159490
rect 329974 159430 330124 159490
rect 330710 159430 330804 159490
rect 331262 159430 331348 159490
rect 332366 159430 332436 159490
rect 333464 159490 333524 160106
rect 333600 159490 333660 160106
rect 334552 159490 334612 160106
rect 335912 159490 335972 160106
rect 336048 159490 336108 160106
rect 337000 159490 337060 160106
rect 338088 159490 338148 160106
rect 338496 159490 338556 160106
rect 339448 159490 339508 160106
rect 340672 159490 340732 160106
rect 341080 159490 341140 160106
rect 341760 159490 341820 160106
rect 333464 159430 333530 159490
rect 333600 159430 333714 159490
rect 334552 159430 334634 159490
rect 327579 158676 327645 158677
rect 327579 158612 327580 158676
rect 327644 158612 327645 158676
rect 327579 158611 327645 158612
rect 328315 158676 328381 158677
rect 328315 158612 328316 158676
rect 328380 158612 328381 158676
rect 328315 158611 328381 158612
rect 328686 158405 328746 159430
rect 329974 158677 330034 159430
rect 330710 158677 330770 159430
rect 331262 158677 331322 159430
rect 332366 158677 332426 159430
rect 329971 158676 330037 158677
rect 329971 158612 329972 158676
rect 330036 158612 330037 158676
rect 329971 158611 330037 158612
rect 330707 158676 330773 158677
rect 330707 158612 330708 158676
rect 330772 158612 330773 158676
rect 330707 158611 330773 158612
rect 331259 158676 331325 158677
rect 331259 158612 331260 158676
rect 331324 158612 331325 158676
rect 331259 158611 331325 158612
rect 332363 158676 332429 158677
rect 332363 158612 332364 158676
rect 332428 158612 332429 158676
rect 332363 158611 332429 158612
rect 328683 158404 328749 158405
rect 328683 158340 328684 158404
rect 328748 158340 328749 158404
rect 328683 158339 328749 158340
rect 333470 158269 333530 159430
rect 333654 158677 333714 159430
rect 334574 158677 334634 159430
rect 335862 159430 335972 159490
rect 336046 159430 336108 159490
rect 336966 159430 337060 159490
rect 338070 159430 338148 159490
rect 338438 159430 338556 159490
rect 339358 159430 339508 159490
rect 340646 159430 340732 159490
rect 341014 159430 341140 159490
rect 341750 159430 341820 159490
rect 342848 159490 342908 160106
rect 343528 159490 343588 160106
rect 343936 159490 343996 160106
rect 345296 159490 345356 160106
rect 342848 159430 342914 159490
rect 343528 159430 343650 159490
rect 343936 159430 344018 159490
rect 335862 158677 335922 159430
rect 336046 158677 336106 159430
rect 336966 158677 337026 159430
rect 333651 158676 333717 158677
rect 333651 158612 333652 158676
rect 333716 158612 333717 158676
rect 333651 158611 333717 158612
rect 334571 158676 334637 158677
rect 334571 158612 334572 158676
rect 334636 158612 334637 158676
rect 334571 158611 334637 158612
rect 335859 158676 335925 158677
rect 335859 158612 335860 158676
rect 335924 158612 335925 158676
rect 335859 158611 335925 158612
rect 336043 158676 336109 158677
rect 336043 158612 336044 158676
rect 336108 158612 336109 158676
rect 336043 158611 336109 158612
rect 336963 158676 337029 158677
rect 336963 158612 336964 158676
rect 337028 158612 337029 158676
rect 336963 158611 337029 158612
rect 338070 158269 338130 159430
rect 338438 158677 338498 159430
rect 339358 158677 339418 159430
rect 338435 158676 338501 158677
rect 338435 158612 338436 158676
rect 338500 158612 338501 158676
rect 338435 158611 338501 158612
rect 339355 158676 339421 158677
rect 339355 158612 339356 158676
rect 339420 158612 339421 158676
rect 339355 158611 339421 158612
rect 333467 158268 333533 158269
rect 333467 158204 333468 158268
rect 333532 158204 333533 158268
rect 333467 158203 333533 158204
rect 338067 158268 338133 158269
rect 338067 158204 338068 158268
rect 338132 158204 338133 158268
rect 338067 158203 338133 158204
rect 326475 158132 326541 158133
rect 326475 158068 326476 158132
rect 326540 158068 326541 158132
rect 326475 158067 326541 158068
rect 325371 157452 325437 157453
rect 325371 157388 325372 157452
rect 325436 157388 325437 157452
rect 325371 157387 325437 157388
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 147454 326414 158000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 151954 330914 158000
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 156454 335414 158000
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 124954 339914 158000
rect 340646 157861 340706 159430
rect 341014 158677 341074 159430
rect 341011 158676 341077 158677
rect 341011 158612 341012 158676
rect 341076 158612 341077 158676
rect 341011 158611 341077 158612
rect 341750 157997 341810 159430
rect 341747 157996 341813 157997
rect 341747 157932 341748 157996
rect 341812 157932 341813 157996
rect 341747 157931 341813 157932
rect 342854 157861 342914 159430
rect 343590 158677 343650 159430
rect 343587 158676 343653 158677
rect 343587 158612 343588 158676
rect 343652 158612 343653 158676
rect 343587 158611 343653 158612
rect 343958 158269 344018 159430
rect 345246 159430 345356 159490
rect 345976 159490 346036 160106
rect 346384 159490 346444 160106
rect 345976 159430 346042 159490
rect 343955 158268 344021 158269
rect 343955 158204 343956 158268
rect 344020 158204 344021 158268
rect 343955 158203 344021 158204
rect 340643 157860 340709 157861
rect 340643 157796 340644 157860
rect 340708 157796 340709 157860
rect 340643 157795 340709 157796
rect 342851 157860 342917 157861
rect 342851 157796 342852 157860
rect 342916 157796 342917 157860
rect 342851 157795 342917 157796
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 129454 344414 158000
rect 345246 157997 345306 159430
rect 345243 157996 345309 157997
rect 345243 157932 345244 157996
rect 345308 157932 345309 157996
rect 345243 157931 345309 157932
rect 345982 157453 346042 159430
rect 346350 159430 346444 159490
rect 347608 159490 347668 160106
rect 348288 159901 348348 160106
rect 348285 159900 348351 159901
rect 348285 159836 348286 159900
rect 348350 159836 348351 159900
rect 348285 159835 348351 159836
rect 348696 159490 348756 160106
rect 349784 159490 349844 160106
rect 351008 159901 351068 160106
rect 351005 159900 351071 159901
rect 351005 159836 351006 159900
rect 351070 159836 351071 159900
rect 351005 159835 351071 159836
rect 351144 159490 351204 160106
rect 347608 159430 347698 159490
rect 348696 159430 348802 159490
rect 349784 159430 349906 159490
rect 346350 157997 346410 159430
rect 347638 158677 347698 159430
rect 347635 158676 347701 158677
rect 347635 158612 347636 158676
rect 347700 158612 347701 158676
rect 347635 158611 347701 158612
rect 348742 158269 348802 159430
rect 348739 158268 348805 158269
rect 348739 158204 348740 158268
rect 348804 158204 348805 158268
rect 348739 158203 348805 158204
rect 346347 157996 346413 157997
rect 346347 157932 346348 157996
rect 346412 157932 346413 157996
rect 346347 157931 346413 157932
rect 345979 157452 346045 157453
rect 345979 157388 345980 157452
rect 346044 157388 346045 157452
rect 345979 157387 346045 157388
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 133954 348914 158000
rect 349846 157453 349906 159430
rect 351134 159430 351204 159490
rect 352232 159490 352292 160106
rect 353320 159490 353380 160106
rect 353592 159629 353652 160106
rect 353589 159628 353655 159629
rect 353589 159564 353590 159628
rect 353654 159564 353655 159628
rect 353589 159563 353655 159564
rect 354408 159490 354468 160106
rect 355768 159490 355828 160106
rect 356040 159901 356100 160106
rect 356037 159900 356103 159901
rect 356037 159836 356038 159900
rect 356102 159836 356103 159900
rect 356037 159835 356103 159836
rect 352232 159430 352298 159490
rect 353320 159430 353402 159490
rect 354408 159430 354506 159490
rect 351134 157453 351194 159430
rect 352238 157453 352298 159430
rect 353342 158269 353402 159430
rect 354446 158677 354506 159430
rect 355734 159430 355828 159490
rect 356992 159490 357052 160106
rect 358080 159490 358140 160106
rect 358488 159901 358548 160106
rect 358485 159900 358551 159901
rect 358485 159836 358486 159900
rect 358550 159836 358551 159900
rect 358485 159835 358551 159836
rect 359168 159490 359228 160106
rect 360936 159901 360996 160106
rect 360933 159900 360999 159901
rect 360933 159836 360934 159900
rect 360998 159836 360999 159900
rect 360933 159835 360999 159836
rect 363520 159490 363580 160106
rect 365968 159629 366028 160106
rect 368280 159901 368340 160106
rect 368277 159900 368343 159901
rect 368277 159836 368278 159900
rect 368342 159836 368343 159900
rect 368277 159835 368343 159836
rect 365965 159628 366031 159629
rect 365965 159564 365966 159628
rect 366030 159564 366031 159628
rect 365965 159563 366031 159564
rect 356992 159430 357082 159490
rect 358080 159430 358186 159490
rect 359168 159430 359290 159490
rect 355734 158677 355794 159430
rect 357022 158677 357082 159430
rect 354443 158676 354509 158677
rect 354443 158612 354444 158676
rect 354508 158612 354509 158676
rect 354443 158611 354509 158612
rect 355731 158676 355797 158677
rect 355731 158612 355732 158676
rect 355796 158612 355797 158676
rect 355731 158611 355797 158612
rect 357019 158676 357085 158677
rect 357019 158612 357020 158676
rect 357084 158612 357085 158676
rect 357019 158611 357085 158612
rect 358126 158541 358186 159430
rect 358123 158540 358189 158541
rect 358123 158476 358124 158540
rect 358188 158476 358189 158540
rect 358123 158475 358189 158476
rect 353339 158268 353405 158269
rect 353339 158204 353340 158268
rect 353404 158204 353405 158268
rect 353339 158203 353405 158204
rect 349843 157452 349909 157453
rect 349843 157388 349844 157452
rect 349908 157388 349909 157452
rect 349843 157387 349909 157388
rect 351131 157452 351197 157453
rect 351131 157388 351132 157452
rect 351196 157388 351197 157452
rect 351131 157387 351197 157388
rect 352235 157452 352301 157453
rect 352235 157388 352236 157452
rect 352300 157388 352301 157452
rect 352235 157387 352301 157388
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 138454 353414 158000
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 142954 357914 158000
rect 359230 157589 359290 159430
rect 363462 159430 363580 159490
rect 371000 159490 371060 160106
rect 373448 159490 373508 160106
rect 371000 159430 371066 159490
rect 363462 158677 363522 159430
rect 371006 158677 371066 159430
rect 373398 159430 373508 159490
rect 375896 159490 375956 160106
rect 378480 159490 378540 160106
rect 380928 159490 380988 160106
rect 383512 159490 383572 160106
rect 385960 159490 386020 160106
rect 388544 159490 388604 160106
rect 375896 159430 376034 159490
rect 378480 159430 378610 159490
rect 380928 159430 381002 159490
rect 383512 159430 383578 159490
rect 373398 158677 373458 159430
rect 375974 158677 376034 159430
rect 378550 158677 378610 159430
rect 380942 158677 381002 159430
rect 383518 158677 383578 159430
rect 385910 159430 386020 159490
rect 388486 159430 388604 159490
rect 390992 159490 391052 160106
rect 393440 159490 393500 160106
rect 395888 159490 395948 160106
rect 398472 159490 398532 160106
rect 390992 159430 391122 159490
rect 393440 159430 393514 159490
rect 385910 158677 385970 159430
rect 388486 158677 388546 159430
rect 391062 158677 391122 159430
rect 393454 158677 393514 159430
rect 395846 159430 395948 159490
rect 398422 159430 398532 159490
rect 400920 159490 400980 160106
rect 403368 159490 403428 160106
rect 405952 159490 406012 160106
rect 400920 159430 401058 159490
rect 403368 159430 403450 159490
rect 405952 159430 406026 159490
rect 395846 158677 395906 159430
rect 398422 158677 398482 159430
rect 400998 158677 401058 159430
rect 403390 158677 403450 159430
rect 405966 158677 406026 159430
rect 363459 158676 363525 158677
rect 363459 158612 363460 158676
rect 363524 158612 363525 158676
rect 363459 158611 363525 158612
rect 371003 158676 371069 158677
rect 371003 158612 371004 158676
rect 371068 158612 371069 158676
rect 371003 158611 371069 158612
rect 373395 158676 373461 158677
rect 373395 158612 373396 158676
rect 373460 158612 373461 158676
rect 373395 158611 373461 158612
rect 375971 158676 376037 158677
rect 375971 158612 375972 158676
rect 376036 158612 376037 158676
rect 375971 158611 376037 158612
rect 378547 158676 378613 158677
rect 378547 158612 378548 158676
rect 378612 158612 378613 158676
rect 378547 158611 378613 158612
rect 380939 158676 381005 158677
rect 380939 158612 380940 158676
rect 381004 158612 381005 158676
rect 380939 158611 381005 158612
rect 383515 158676 383581 158677
rect 383515 158612 383516 158676
rect 383580 158612 383581 158676
rect 383515 158611 383581 158612
rect 385907 158676 385973 158677
rect 385907 158612 385908 158676
rect 385972 158612 385973 158676
rect 385907 158611 385973 158612
rect 388483 158676 388549 158677
rect 388483 158612 388484 158676
rect 388548 158612 388549 158676
rect 388483 158611 388549 158612
rect 391059 158676 391125 158677
rect 391059 158612 391060 158676
rect 391124 158612 391125 158676
rect 391059 158611 391125 158612
rect 393451 158676 393517 158677
rect 393451 158612 393452 158676
rect 393516 158612 393517 158676
rect 393451 158611 393517 158612
rect 395843 158676 395909 158677
rect 395843 158612 395844 158676
rect 395908 158612 395909 158676
rect 395843 158611 395909 158612
rect 398419 158676 398485 158677
rect 398419 158612 398420 158676
rect 398484 158612 398485 158676
rect 398419 158611 398485 158612
rect 400995 158676 401061 158677
rect 400995 158612 400996 158676
rect 401060 158612 401061 158676
rect 400995 158611 401061 158612
rect 403387 158676 403453 158677
rect 403387 158612 403388 158676
rect 403452 158612 403453 158676
rect 403387 158611 403453 158612
rect 405963 158676 406029 158677
rect 405963 158612 405964 158676
rect 406028 158612 406029 158676
rect 405963 158611 406029 158612
rect 359227 157588 359293 157589
rect 359227 157524 359228 157588
rect 359292 157524 359293 157588
rect 359227 157523 359293 157524
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 147454 362414 158000
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 151954 366914 158000
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 156454 371414 158000
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 124954 375914 158000
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 129454 380414 158000
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 133954 384914 158000
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 138454 389414 158000
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 142954 393914 158000
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 147454 398414 158000
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 151954 402914 158000
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 156454 407414 158000
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 124954 411914 158000
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 129454 416414 158000
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 133954 420914 158000
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 138454 425414 158000
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 142954 429914 158000
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 147454 434414 158000
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 437430 3501 437490 287675
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 437611 247620 437677 247621
rect 437611 247556 437612 247620
rect 437676 247556 437677 247620
rect 437611 247555 437677 247556
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 437427 3500 437493 3501
rect 437427 3436 437428 3500
rect 437492 3436 437493 3500
rect 437427 3435 437493 3436
rect 437614 3365 437674 247555
rect 437795 245308 437861 245309
rect 438294 245308 438914 259398
rect 437795 245244 437796 245308
rect 437860 245244 437861 245308
rect 437795 245243 437861 245244
rect 437798 3637 437858 245243
rect 438294 151954 438914 158000
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 437795 3636 437861 3637
rect 437795 3572 437796 3636
rect 437860 3572 437861 3636
rect 437795 3571 437861 3572
rect 437611 3364 437677 3365
rect 437611 3300 437612 3364
rect 437676 3300 437677 3364
rect 437611 3299 437677 3300
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 -1306 438914 7398
rect 439086 3501 439146 298691
rect 439454 4045 439514 302907
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 439451 4044 439517 4045
rect 439451 3980 439452 4044
rect 439516 3980 439517 4044
rect 439451 3979 439517 3980
rect 439083 3500 439149 3501
rect 439083 3436 439084 3500
rect 439148 3436 439149 3500
rect 439083 3435 439149 3436
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 220328 547718 220564 547954
rect 220328 547398 220564 547634
rect 356056 547718 356292 547954
rect 356056 547398 356292 547634
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 220328 511718 220564 511954
rect 220328 511398 220564 511634
rect 356056 511718 356292 511954
rect 356056 511398 356292 511634
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 249610 439718 249846 439954
rect 249610 439398 249846 439634
rect 280330 439718 280566 439954
rect 280330 439398 280566 439634
rect 311050 439718 311286 439954
rect 311050 439398 311286 439634
rect 341770 439718 342006 439954
rect 341770 439398 342006 439634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 234250 435218 234486 435454
rect 234250 434898 234486 435134
rect 264970 435218 265206 435454
rect 264970 434898 265206 435134
rect 295690 435218 295926 435454
rect 295690 434898 295926 435134
rect 326410 435218 326646 435454
rect 326410 434898 326646 435134
rect 357130 435218 357366 435454
rect 357130 434898 357366 435134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 249610 403718 249846 403954
rect 249610 403398 249846 403634
rect 280330 403718 280566 403954
rect 280330 403398 280566 403634
rect 311050 403718 311286 403954
rect 311050 403398 311286 403634
rect 341770 403718 342006 403954
rect 341770 403398 342006 403634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 234250 399218 234486 399454
rect 234250 398898 234486 399134
rect 264970 399218 265206 399454
rect 264970 398898 265206 399134
rect 295690 399218 295926 399454
rect 295690 398898 295926 399134
rect 326410 399218 326646 399454
rect 326410 398898 326646 399134
rect 357130 399218 357366 399454
rect 357130 398898 357366 399134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 249610 367718 249846 367954
rect 249610 367398 249846 367634
rect 280330 367718 280566 367954
rect 280330 367398 280566 367634
rect 311050 367718 311286 367954
rect 311050 367398 311286 367634
rect 341770 367718 342006 367954
rect 341770 367398 342006 367634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 234250 363218 234486 363454
rect 234250 362898 234486 363134
rect 264970 363218 265206 363454
rect 264970 362898 265206 363134
rect 295690 363218 295926 363454
rect 295690 362898 295926 363134
rect 326410 363218 326646 363454
rect 326410 362898 326646 363134
rect 357130 363218 357366 363454
rect 357130 362898 357366 363134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 249610 331718 249846 331954
rect 249610 331398 249846 331634
rect 280330 331718 280566 331954
rect 280330 331398 280566 331634
rect 311050 331718 311286 331954
rect 311050 331398 311286 331634
rect 341770 331718 342006 331954
rect 341770 331398 342006 331634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 234250 327218 234486 327454
rect 234250 326898 234486 327134
rect 264970 327218 265206 327454
rect 264970 326898 265206 327134
rect 295690 327218 295926 327454
rect 295690 326898 295926 327134
rect 326410 327218 326646 327454
rect 326410 326898 326646 327134
rect 357130 327218 357366 327454
rect 357130 326898 357366 327134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 100328 223718 100564 223954
rect 100328 223398 100564 223634
rect 236056 223718 236292 223954
rect 236056 223398 236292 223634
rect 101008 219218 101244 219454
rect 101008 218898 101244 219134
rect 235376 219218 235612 219454
rect 235376 218898 235612 219134
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 100328 187718 100564 187954
rect 100328 187398 100564 187634
rect 236056 187718 236292 187954
rect 236056 187398 236292 187634
rect 101008 183218 101244 183454
rect 101008 182898 101244 183134
rect 235376 183218 235612 183454
rect 235376 182898 235612 183134
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 300328 223718 300564 223954
rect 300328 223398 300564 223634
rect 436056 223718 436292 223954
rect 436056 223398 436292 223634
rect 301008 219218 301244 219454
rect 301008 218898 301244 219134
rect 435376 219218 435612 219454
rect 435376 218898 435612 219134
rect 300328 187718 300564 187954
rect 300328 187398 300564 187634
rect 436056 187718 436292 187954
rect 436056 187398 436292 187634
rect 301008 183218 301244 183454
rect 301008 182898 301244 183134
rect 435376 183218 435612 183454
rect 435376 182898 435612 183134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 220328 547954
rect 220564 547718 356056 547954
rect 356292 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 220328 547634
rect 220564 547398 356056 547634
rect 356292 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 220328 511954
rect 220564 511718 356056 511954
rect 356292 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 220328 511634
rect 220564 511398 356056 511634
rect 356292 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 249610 439954
rect 249846 439718 280330 439954
rect 280566 439718 311050 439954
rect 311286 439718 341770 439954
rect 342006 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 249610 439634
rect 249846 439398 280330 439634
rect 280566 439398 311050 439634
rect 311286 439398 341770 439634
rect 342006 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 234250 435454
rect 234486 435218 264970 435454
rect 265206 435218 295690 435454
rect 295926 435218 326410 435454
rect 326646 435218 357130 435454
rect 357366 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 234250 435134
rect 234486 434898 264970 435134
rect 265206 434898 295690 435134
rect 295926 434898 326410 435134
rect 326646 434898 357130 435134
rect 357366 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 249610 403954
rect 249846 403718 280330 403954
rect 280566 403718 311050 403954
rect 311286 403718 341770 403954
rect 342006 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 249610 403634
rect 249846 403398 280330 403634
rect 280566 403398 311050 403634
rect 311286 403398 341770 403634
rect 342006 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 234250 399454
rect 234486 399218 264970 399454
rect 265206 399218 295690 399454
rect 295926 399218 326410 399454
rect 326646 399218 357130 399454
rect 357366 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 234250 399134
rect 234486 398898 264970 399134
rect 265206 398898 295690 399134
rect 295926 398898 326410 399134
rect 326646 398898 357130 399134
rect 357366 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 249610 367954
rect 249846 367718 280330 367954
rect 280566 367718 311050 367954
rect 311286 367718 341770 367954
rect 342006 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 249610 367634
rect 249846 367398 280330 367634
rect 280566 367398 311050 367634
rect 311286 367398 341770 367634
rect 342006 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 234250 363454
rect 234486 363218 264970 363454
rect 265206 363218 295690 363454
rect 295926 363218 326410 363454
rect 326646 363218 357130 363454
rect 357366 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 234250 363134
rect 234486 362898 264970 363134
rect 265206 362898 295690 363134
rect 295926 362898 326410 363134
rect 326646 362898 357130 363134
rect 357366 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 249610 331954
rect 249846 331718 280330 331954
rect 280566 331718 311050 331954
rect 311286 331718 341770 331954
rect 342006 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 249610 331634
rect 249846 331398 280330 331634
rect 280566 331398 311050 331634
rect 311286 331398 341770 331634
rect 342006 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 234250 327454
rect 234486 327218 264970 327454
rect 265206 327218 295690 327454
rect 295926 327218 326410 327454
rect 326646 327218 357130 327454
rect 357366 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 234250 327134
rect 234486 326898 264970 327134
rect 265206 326898 295690 327134
rect 295926 326898 326410 327134
rect 326646 326898 357130 327134
rect 357366 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 100328 223954
rect 100564 223718 236056 223954
rect 236292 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 300328 223954
rect 300564 223718 436056 223954
rect 436292 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 100328 223634
rect 100564 223398 236056 223634
rect 236292 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 300328 223634
rect 300564 223398 436056 223634
rect 436292 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 101008 219454
rect 101244 219218 235376 219454
rect 235612 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 301008 219454
rect 301244 219218 435376 219454
rect 435612 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 101008 219134
rect 101244 218898 235376 219134
rect 235612 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 301008 219134
rect 301244 218898 435376 219134
rect 435612 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 100328 187954
rect 100564 187718 236056 187954
rect 236292 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 300328 187954
rect 300564 187718 436056 187954
rect 436292 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 100328 187634
rect 100564 187398 236056 187634
rect 236292 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 300328 187634
rect 300564 187398 436056 187634
rect 436292 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 101008 183454
rect 101244 183218 235376 183454
rect 235612 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 301008 183454
rect 301244 183218 435376 183454
rect 435612 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 101008 183134
rect 101244 182898 235376 183134
rect 235612 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 301008 183134
rect 301244 182898 435376 183134
rect 435612 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  dram_inst
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst_A
timestamp 0
transform 1 0 100000 0 1 160000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst_B
timestamp 0
transform 1 0 300000 0 1 160000
box 0 0 136620 83308
use rvj1_caravel_soc  rvj1_soc
timestamp 0
transform 1 0 230000 0 1 310400
box 14 0 130994 133208
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 245308 110414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 245308 146414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 245308 182414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 245308 218414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 565308 218414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 565308 254414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 565308 290414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 245308 326414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 565308 326414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 245308 362414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 445608 362414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 245308 398414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 245308 434414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7654 11414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7654 47414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7654 83414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7654 119414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 245308 119414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7654 155414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 245308 155414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7654 191414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 245308 191414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7654 227414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 245308 227414 478000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 565308 227414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7654 263414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 565308 263414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7654 299414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 245308 299414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 565308 299414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7654 335414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 245308 335414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 565308 335414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7654 371414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 245308 371414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7654 407414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 245308 407414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7654 443414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7654 479414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7654 515414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7654 551414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 11866 592650 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 47866 592650 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 83866 592650 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 119866 592650 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 155866 592650 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 191866 592650 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 227866 592650 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 263866 592650 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 299866 592650 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 335866 592650 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 371866 592650 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 407866 592650 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 443866 592650 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 479866 592650 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 515866 592650 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 551866 592650 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 587866 592650 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 623866 592650 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 659866 592650 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 695866 592650 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 19794 -7654 20414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 55794 -7654 56414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 127794 -7654 128414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 127794 245308 128414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 163794 -7654 164414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 163794 245308 164414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 199794 -7654 200414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 199794 245308 200414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 -7654 236414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 565308 236414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 565308 272414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 -7654 308414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 565308 308414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 -7654 344414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 565308 344414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 379794 -7654 380414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 379794 245308 380414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 415794 -7654 416414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 415794 245308 416414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 487794 -7654 488414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 523794 -7654 524414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 559794 -7654 560414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 20866 592650 21486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 56866 592650 57486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 128866 592650 129486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 164866 592650 165486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 200866 592650 201486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 236866 592650 237486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 308866 592650 309486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 344866 592650 345486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 380866 592650 381486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 416866 592650 417486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 488866 592650 489486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 524866 592650 525486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 560866 592650 561486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 596866 592650 597486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 668866 592650 669486 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 28794 -7654 29414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 64794 -7654 65414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 100794 -7654 101414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 100794 245308 101414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 136794 -7654 137414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 136794 245308 137414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 172794 -7654 173414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 172794 245308 173414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 208794 -7654 209414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 208794 245308 209414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 -7654 245414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 565308 245414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 -7654 281414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 565308 281414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 -7654 317414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 245308 317414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 565308 317414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 -7654 353414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 245308 353414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 565308 353414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 388794 -7654 389414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 388794 245308 389414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 424794 -7654 425414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 424794 245308 425414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 460794 -7654 461414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 496794 -7654 497414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 532794 -7654 533414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 568794 -7654 569414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 29866 592650 30486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 65866 592650 66486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 101866 592650 102486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 137866 592650 138486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 173866 592650 174486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 209866 592650 210486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 245866 592650 246486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 281866 592650 282486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 317866 592650 318486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 353866 592650 354486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 389866 592650 390486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 425866 592650 426486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 461866 592650 462486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 497866 592650 498486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 533866 592650 534486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 569866 592650 570486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 605866 592650 606486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 641866 592650 642486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 677866 592650 678486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 24294 -7654 24914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 60294 -7654 60914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 96294 -7654 96914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 132294 -7654 132914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 132294 245308 132914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 168294 -7654 168914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 168294 245308 168914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 204294 -7654 204914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 204294 245308 204914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 -7654 240914 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 565308 240914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 -7654 276914 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 565308 276914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 -7654 312914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 565308 312914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 -7654 348914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 565308 348914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 384294 -7654 384914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 384294 245308 384914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 420294 -7654 420914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 420294 245308 420914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 456294 -7654 456914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 492294 -7654 492914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 528294 -7654 528914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 564294 -7654 564914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 25366 592650 25986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 61366 592650 61986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 97366 592650 97986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 133366 592650 133986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 169366 592650 169986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 205366 592650 205986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 241366 592650 241986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 277366 592650 277986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 313366 592650 313986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 349366 592650 349986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 385366 592650 385986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 421366 592650 421986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 457366 592650 457986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 493366 592650 493986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 529366 592650 529986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 565366 592650 565986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 601366 592650 601986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 637366 592650 637986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 673366 592650 673986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7654 33914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7654 69914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7654 105914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 245308 105914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7654 141914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 245308 141914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7654 177914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 245308 177914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7654 213914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 245308 213914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7654 249914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 565308 249914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7654 285914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 565308 285914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7654 321914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 245308 321914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 565308 321914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7654 357914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 245308 357914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 565308 357914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7654 393914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 245308 393914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7654 429914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 245308 429914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7654 465914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7654 501914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7654 537914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7654 573914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 34366 592650 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 70366 592650 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 106366 592650 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 142366 592650 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 178366 592650 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 214366 592650 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 250366 592650 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 286366 592650 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 322366 592650 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 358366 592650 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 394366 592650 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 430366 592650 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 466366 592650 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 502366 592650 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 538366 592650 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 574366 592650 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 610366 592650 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 646366 592650 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 682366 592650 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7654 6914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7654 42914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7654 78914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7654 114914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 245308 114914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7654 150914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 245308 150914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7654 186914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 245308 186914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7654 222914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 245308 222914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 565308 222914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7654 258914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 565308 258914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7654 294914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 565308 294914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7654 330914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 245308 330914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 565308 330914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7654 366914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 245308 366914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7654 402914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 245308 402914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7654 438914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 245308 438914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7654 474914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7654 510914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7654 546914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7654 582914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 7366 592650 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 43366 592650 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 79366 592650 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 115366 592650 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 151366 592650 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 187366 592650 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 223366 592650 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 259366 592650 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 295366 592650 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 331366 592650 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 367366 592650 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 403366 592650 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 439366 592650 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 475366 592650 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 511366 592650 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 547366 592650 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 583366 592650 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 619366 592650 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 655366 592650 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 691366 592650 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 15294 -7654 15914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 51294 -7654 51914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 87294 -7654 87914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 123294 -7654 123914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 123294 245308 123914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 159294 -7654 159914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 159294 245308 159914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 195294 -7654 195914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 195294 245308 195914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 -7654 231914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 245308 231914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 565308 231914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 -7654 267914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 565308 267914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 -7654 303914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 245308 303914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 565308 303914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 -7654 339914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 245308 339914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 565308 339914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 375294 -7654 375914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 375294 245308 375914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 411294 -7654 411914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 411294 245308 411914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 447294 -7654 447914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 483294 -7654 483914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 519294 -7654 519914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 555294 -7654 555914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 16366 592650 16986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 52366 592650 52986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 88366 592650 88986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 124366 592650 124986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 160366 592650 160986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 196366 592650 196986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 232366 592650 232986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 268366 592650 268986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 304366 592650 304986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 340366 592650 340986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 376366 592650 376986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 412366 592650 412986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 448366 592650 448986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 484366 592650 484986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 520366 592650 520986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 556366 592650 556986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 592366 592650 592986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 628366 592650 628986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 664366 592650 664986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 700366 592650 700986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
