magic
tech sky130A
magscale 1 2
timestamp 1654694221
<< obsli1 >>
rect 1104 2159 129904 130577
<< obsm1 >>
rect 14 212 130994 131708
<< metal2 >>
rect 386 132408 442 133208
rect 1122 132408 1178 133208
rect 1858 132408 1914 133208
rect 2686 132408 2742 133208
rect 3422 132408 3478 133208
rect 4250 132408 4306 133208
rect 4986 132408 5042 133208
rect 5814 132408 5870 133208
rect 6550 132408 6606 133208
rect 7286 132408 7342 133208
rect 8114 132408 8170 133208
rect 8850 132408 8906 133208
rect 9678 132408 9734 133208
rect 10414 132408 10470 133208
rect 11242 132408 11298 133208
rect 11978 132408 12034 133208
rect 12714 132408 12770 133208
rect 13542 132408 13598 133208
rect 14278 132408 14334 133208
rect 15106 132408 15162 133208
rect 15842 132408 15898 133208
rect 16670 132408 16726 133208
rect 17406 132408 17462 133208
rect 18142 132408 18198 133208
rect 18970 132408 19026 133208
rect 19706 132408 19762 133208
rect 20534 132408 20590 133208
rect 21270 132408 21326 133208
rect 22098 132408 22154 133208
rect 22834 132408 22890 133208
rect 23570 132408 23626 133208
rect 24398 132408 24454 133208
rect 25134 132408 25190 133208
rect 25962 132408 26018 133208
rect 26698 132408 26754 133208
rect 27526 132408 27582 133208
rect 28262 132408 28318 133208
rect 28998 132408 29054 133208
rect 29826 132408 29882 133208
rect 30562 132408 30618 133208
rect 31390 132408 31446 133208
rect 32126 132408 32182 133208
rect 32954 132408 33010 133208
rect 33690 132408 33746 133208
rect 34518 132408 34574 133208
rect 35254 132408 35310 133208
rect 35990 132408 36046 133208
rect 36818 132408 36874 133208
rect 37554 132408 37610 133208
rect 38382 132408 38438 133208
rect 39118 132408 39174 133208
rect 39946 132408 40002 133208
rect 40682 132408 40738 133208
rect 41418 132408 41474 133208
rect 42246 132408 42302 133208
rect 42982 132408 43038 133208
rect 43810 132408 43866 133208
rect 44546 132408 44602 133208
rect 45374 132408 45430 133208
rect 46110 132408 46166 133208
rect 46846 132408 46902 133208
rect 47674 132408 47730 133208
rect 48410 132408 48466 133208
rect 49238 132408 49294 133208
rect 49974 132408 50030 133208
rect 50802 132408 50858 133208
rect 51538 132408 51594 133208
rect 52274 132408 52330 133208
rect 53102 132408 53158 133208
rect 53838 132408 53894 133208
rect 54666 132408 54722 133208
rect 55402 132408 55458 133208
rect 56230 132408 56286 133208
rect 56966 132408 57022 133208
rect 57702 132408 57758 133208
rect 58530 132408 58586 133208
rect 59266 132408 59322 133208
rect 60094 132408 60150 133208
rect 60830 132408 60886 133208
rect 61658 132408 61714 133208
rect 62394 132408 62450 133208
rect 63130 132408 63186 133208
rect 63958 132408 64014 133208
rect 64694 132408 64750 133208
rect 65522 132408 65578 133208
rect 66258 132408 66314 133208
rect 67086 132408 67142 133208
rect 67822 132408 67878 133208
rect 68650 132408 68706 133208
rect 69386 132408 69442 133208
rect 70122 132408 70178 133208
rect 70950 132408 71006 133208
rect 71686 132408 71742 133208
rect 72514 132408 72570 133208
rect 73250 132408 73306 133208
rect 74078 132408 74134 133208
rect 74814 132408 74870 133208
rect 75550 132408 75606 133208
rect 76378 132408 76434 133208
rect 77114 132408 77170 133208
rect 77942 132408 77998 133208
rect 78678 132408 78734 133208
rect 79506 132408 79562 133208
rect 80242 132408 80298 133208
rect 80978 132408 81034 133208
rect 81806 132408 81862 133208
rect 82542 132408 82598 133208
rect 83370 132408 83426 133208
rect 84106 132408 84162 133208
rect 84934 132408 84990 133208
rect 85670 132408 85726 133208
rect 86406 132408 86462 133208
rect 87234 132408 87290 133208
rect 87970 132408 88026 133208
rect 88798 132408 88854 133208
rect 89534 132408 89590 133208
rect 90362 132408 90418 133208
rect 91098 132408 91154 133208
rect 91834 132408 91890 133208
rect 92662 132408 92718 133208
rect 93398 132408 93454 133208
rect 94226 132408 94282 133208
rect 94962 132408 95018 133208
rect 95790 132408 95846 133208
rect 96526 132408 96582 133208
rect 97262 132408 97318 133208
rect 98090 132408 98146 133208
rect 98826 132408 98882 133208
rect 99654 132408 99710 133208
rect 100390 132408 100446 133208
rect 101218 132408 101274 133208
rect 101954 132408 102010 133208
rect 102782 132408 102838 133208
rect 103518 132408 103574 133208
rect 104254 132408 104310 133208
rect 105082 132408 105138 133208
rect 105818 132408 105874 133208
rect 106646 132408 106702 133208
rect 107382 132408 107438 133208
rect 108210 132408 108266 133208
rect 108946 132408 109002 133208
rect 109682 132408 109738 133208
rect 110510 132408 110566 133208
rect 111246 132408 111302 133208
rect 112074 132408 112130 133208
rect 112810 132408 112866 133208
rect 113638 132408 113694 133208
rect 114374 132408 114430 133208
rect 115110 132408 115166 133208
rect 115938 132408 115994 133208
rect 116674 132408 116730 133208
rect 117502 132408 117558 133208
rect 118238 132408 118294 133208
rect 119066 132408 119122 133208
rect 119802 132408 119858 133208
rect 120538 132408 120594 133208
rect 121366 132408 121422 133208
rect 122102 132408 122158 133208
rect 122930 132408 122986 133208
rect 123666 132408 123722 133208
rect 124494 132408 124550 133208
rect 125230 132408 125286 133208
rect 125966 132408 126022 133208
rect 126794 132408 126850 133208
rect 127530 132408 127586 133208
rect 128358 132408 128414 133208
rect 129094 132408 129150 133208
rect 129922 132408 129978 133208
rect 130658 132408 130714 133208
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 754 0 810 800
rect 938 0 994 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10690 0 10746 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19890 0 19946 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64234 0 64290 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68098 0 68154 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 69018 0 69074 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72698 0 72754 800
rect 72882 0 72938 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 73986 0 74042 800
rect 74170 0 74226 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76838 0 76894 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78586 0 78642 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79230 0 79286 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82266 0 82322 800
rect 82450 0 82506 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83554 0 83610 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86130 0 86186 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86774 0 86830 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89442 0 89498 800
rect 89626 0 89682 800
rect 89810 0 89866 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91834 0 91890 800
rect 92018 0 92074 800
rect 92202 0 92258 800
rect 92478 0 92534 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95054 0 95110 800
rect 95330 0 95386 800
rect 95514 0 95570 800
rect 95698 0 95754 800
rect 95974 0 96030 800
rect 96158 0 96214 800
rect 96342 0 96398 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 97906 0 97962 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98550 0 98606 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99194 0 99250 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100298 0 100354 800
rect 100482 0 100538 800
rect 100758 0 100814 800
rect 100942 0 100998 800
rect 101126 0 101182 800
rect 101402 0 101458 800
rect 101586 0 101642 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102690 0 102746 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103334 0 103390 800
rect 103518 0 103574 800
rect 103794 0 103850 800
rect 103978 0 104034 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104622 0 104678 800
rect 104898 0 104954 800
rect 105082 0 105138 800
rect 105266 0 105322 800
rect 105542 0 105598 800
rect 105726 0 105782 800
rect 105910 0 105966 800
rect 106186 0 106242 800
rect 106370 0 106426 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107474 0 107530 800
rect 107658 0 107714 800
rect 107934 0 107990 800
rect 108118 0 108174 800
rect 108302 0 108358 800
rect 108578 0 108634 800
rect 108762 0 108818 800
rect 108946 0 109002 800
rect 109222 0 109278 800
rect 109406 0 109462 800
rect 109682 0 109738 800
rect 109866 0 109922 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110510 0 110566 800
rect 110694 0 110750 800
rect 110970 0 111026 800
rect 111154 0 111210 800
rect 111338 0 111394 800
rect 111614 0 111670 800
rect 111798 0 111854 800
rect 112074 0 112130 800
rect 112258 0 112314 800
rect 112442 0 112498 800
rect 112718 0 112774 800
rect 112902 0 112958 800
rect 113086 0 113142 800
rect 113362 0 113418 800
rect 113546 0 113602 800
rect 113730 0 113786 800
rect 114006 0 114062 800
rect 114190 0 114246 800
rect 114466 0 114522 800
rect 114650 0 114706 800
rect 114834 0 114890 800
rect 115110 0 115166 800
rect 115294 0 115350 800
rect 115478 0 115534 800
rect 115754 0 115810 800
rect 115938 0 115994 800
rect 116122 0 116178 800
rect 116398 0 116454 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117042 0 117098 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117686 0 117742 800
rect 117870 0 117926 800
rect 118146 0 118202 800
rect 118330 0 118386 800
rect 118514 0 118570 800
rect 118790 0 118846 800
rect 118974 0 119030 800
rect 119250 0 119306 800
rect 119434 0 119490 800
rect 119618 0 119674 800
rect 119894 0 119950 800
rect 120078 0 120134 800
rect 120262 0 120318 800
rect 120538 0 120594 800
rect 120722 0 120778 800
rect 120906 0 120962 800
rect 121182 0 121238 800
rect 121366 0 121422 800
rect 121642 0 121698 800
rect 121826 0 121882 800
rect 122010 0 122066 800
rect 122286 0 122342 800
rect 122470 0 122526 800
rect 122654 0 122710 800
rect 122930 0 122986 800
rect 123114 0 123170 800
rect 123298 0 123354 800
rect 123574 0 123630 800
rect 123758 0 123814 800
rect 124034 0 124090 800
rect 124218 0 124274 800
rect 124402 0 124458 800
rect 124678 0 124734 800
rect 124862 0 124918 800
rect 125046 0 125102 800
rect 125322 0 125378 800
rect 125506 0 125562 800
rect 125690 0 125746 800
rect 125966 0 126022 800
rect 126150 0 126206 800
rect 126426 0 126482 800
rect 126610 0 126666 800
rect 126794 0 126850 800
rect 127070 0 127126 800
rect 127254 0 127310 800
rect 127438 0 127494 800
rect 127714 0 127770 800
rect 127898 0 127954 800
rect 128082 0 128138 800
rect 128358 0 128414 800
rect 128542 0 128598 800
rect 128818 0 128874 800
rect 129002 0 129058 800
rect 129186 0 129242 800
rect 129462 0 129518 800
rect 129646 0 129702 800
rect 129830 0 129886 800
rect 130106 0 130162 800
rect 130290 0 130346 800
rect 130474 0 130530 800
rect 130750 0 130806 800
rect 130934 0 130990 800
<< obsm2 >>
rect 20 132352 330 132546
rect 498 132352 1066 132546
rect 1234 132352 1802 132546
rect 1970 132352 2630 132546
rect 2798 132352 3366 132546
rect 3534 132352 4194 132546
rect 4362 132352 4930 132546
rect 5098 132352 5758 132546
rect 5926 132352 6494 132546
rect 6662 132352 7230 132546
rect 7398 132352 8058 132546
rect 8226 132352 8794 132546
rect 8962 132352 9622 132546
rect 9790 132352 10358 132546
rect 10526 132352 11186 132546
rect 11354 132352 11922 132546
rect 12090 132352 12658 132546
rect 12826 132352 13486 132546
rect 13654 132352 14222 132546
rect 14390 132352 15050 132546
rect 15218 132352 15786 132546
rect 15954 132352 16614 132546
rect 16782 132352 17350 132546
rect 17518 132352 18086 132546
rect 18254 132352 18914 132546
rect 19082 132352 19650 132546
rect 19818 132352 20478 132546
rect 20646 132352 21214 132546
rect 21382 132352 22042 132546
rect 22210 132352 22778 132546
rect 22946 132352 23514 132546
rect 23682 132352 24342 132546
rect 24510 132352 25078 132546
rect 25246 132352 25906 132546
rect 26074 132352 26642 132546
rect 26810 132352 27470 132546
rect 27638 132352 28206 132546
rect 28374 132352 28942 132546
rect 29110 132352 29770 132546
rect 29938 132352 30506 132546
rect 30674 132352 31334 132546
rect 31502 132352 32070 132546
rect 32238 132352 32898 132546
rect 33066 132352 33634 132546
rect 33802 132352 34462 132546
rect 34630 132352 35198 132546
rect 35366 132352 35934 132546
rect 36102 132352 36762 132546
rect 36930 132352 37498 132546
rect 37666 132352 38326 132546
rect 38494 132352 39062 132546
rect 39230 132352 39890 132546
rect 40058 132352 40626 132546
rect 40794 132352 41362 132546
rect 41530 132352 42190 132546
rect 42358 132352 42926 132546
rect 43094 132352 43754 132546
rect 43922 132352 44490 132546
rect 44658 132352 45318 132546
rect 45486 132352 46054 132546
rect 46222 132352 46790 132546
rect 46958 132352 47618 132546
rect 47786 132352 48354 132546
rect 48522 132352 49182 132546
rect 49350 132352 49918 132546
rect 50086 132352 50746 132546
rect 50914 132352 51482 132546
rect 51650 132352 52218 132546
rect 52386 132352 53046 132546
rect 53214 132352 53782 132546
rect 53950 132352 54610 132546
rect 54778 132352 55346 132546
rect 55514 132352 56174 132546
rect 56342 132352 56910 132546
rect 57078 132352 57646 132546
rect 57814 132352 58474 132546
rect 58642 132352 59210 132546
rect 59378 132352 60038 132546
rect 60206 132352 60774 132546
rect 60942 132352 61602 132546
rect 61770 132352 62338 132546
rect 62506 132352 63074 132546
rect 63242 132352 63902 132546
rect 64070 132352 64638 132546
rect 64806 132352 65466 132546
rect 65634 132352 66202 132546
rect 66370 132352 67030 132546
rect 67198 132352 67766 132546
rect 67934 132352 68594 132546
rect 68762 132352 69330 132546
rect 69498 132352 70066 132546
rect 70234 132352 70894 132546
rect 71062 132352 71630 132546
rect 71798 132352 72458 132546
rect 72626 132352 73194 132546
rect 73362 132352 74022 132546
rect 74190 132352 74758 132546
rect 74926 132352 75494 132546
rect 75662 132352 76322 132546
rect 76490 132352 77058 132546
rect 77226 132352 77886 132546
rect 78054 132352 78622 132546
rect 78790 132352 79450 132546
rect 79618 132352 80186 132546
rect 80354 132352 80922 132546
rect 81090 132352 81750 132546
rect 81918 132352 82486 132546
rect 82654 132352 83314 132546
rect 83482 132352 84050 132546
rect 84218 132352 84878 132546
rect 85046 132352 85614 132546
rect 85782 132352 86350 132546
rect 86518 132352 87178 132546
rect 87346 132352 87914 132546
rect 88082 132352 88742 132546
rect 88910 132352 89478 132546
rect 89646 132352 90306 132546
rect 90474 132352 91042 132546
rect 91210 132352 91778 132546
rect 91946 132352 92606 132546
rect 92774 132352 93342 132546
rect 93510 132352 94170 132546
rect 94338 132352 94906 132546
rect 95074 132352 95734 132546
rect 95902 132352 96470 132546
rect 96638 132352 97206 132546
rect 97374 132352 98034 132546
rect 98202 132352 98770 132546
rect 98938 132352 99598 132546
rect 99766 132352 100334 132546
rect 100502 132352 101162 132546
rect 101330 132352 101898 132546
rect 102066 132352 102726 132546
rect 102894 132352 103462 132546
rect 103630 132352 104198 132546
rect 104366 132352 105026 132546
rect 105194 132352 105762 132546
rect 105930 132352 106590 132546
rect 106758 132352 107326 132546
rect 107494 132352 108154 132546
rect 108322 132352 108890 132546
rect 109058 132352 109626 132546
rect 109794 132352 110454 132546
rect 110622 132352 111190 132546
rect 111358 132352 112018 132546
rect 112186 132352 112754 132546
rect 112922 132352 113582 132546
rect 113750 132352 114318 132546
rect 114486 132352 115054 132546
rect 115222 132352 115882 132546
rect 116050 132352 116618 132546
rect 116786 132352 117446 132546
rect 117614 132352 118182 132546
rect 118350 132352 119010 132546
rect 119178 132352 119746 132546
rect 119914 132352 120482 132546
rect 120650 132352 121310 132546
rect 121478 132352 122046 132546
rect 122214 132352 122874 132546
rect 123042 132352 123610 132546
rect 123778 132352 124438 132546
rect 124606 132352 125174 132546
rect 125342 132352 125910 132546
rect 126078 132352 126738 132546
rect 126906 132352 127474 132546
rect 127642 132352 128302 132546
rect 128470 132352 129038 132546
rect 129206 132352 129866 132546
rect 130034 132352 130602 132546
rect 130770 132352 130988 132546
rect 20 856 130988 132352
rect 20 206 54 856
rect 222 206 238 856
rect 406 206 422 856
rect 590 206 698 856
rect 866 206 882 856
rect 1050 206 1066 856
rect 1234 206 1342 856
rect 1510 206 1526 856
rect 1694 206 1710 856
rect 1878 206 1986 856
rect 2154 206 2170 856
rect 2338 206 2354 856
rect 2522 206 2630 856
rect 2798 206 2814 856
rect 2982 206 3090 856
rect 3258 206 3274 856
rect 3442 206 3458 856
rect 3626 206 3734 856
rect 3902 206 3918 856
rect 4086 206 4102 856
rect 4270 206 4378 856
rect 4546 206 4562 856
rect 4730 206 4746 856
rect 4914 206 5022 856
rect 5190 206 5206 856
rect 5374 206 5482 856
rect 5650 206 5666 856
rect 5834 206 5850 856
rect 6018 206 6126 856
rect 6294 206 6310 856
rect 6478 206 6494 856
rect 6662 206 6770 856
rect 6938 206 6954 856
rect 7122 206 7138 856
rect 7306 206 7414 856
rect 7582 206 7598 856
rect 7766 206 7874 856
rect 8042 206 8058 856
rect 8226 206 8242 856
rect 8410 206 8518 856
rect 8686 206 8702 856
rect 8870 206 8886 856
rect 9054 206 9162 856
rect 9330 206 9346 856
rect 9514 206 9530 856
rect 9698 206 9806 856
rect 9974 206 9990 856
rect 10158 206 10266 856
rect 10434 206 10450 856
rect 10618 206 10634 856
rect 10802 206 10910 856
rect 11078 206 11094 856
rect 11262 206 11278 856
rect 11446 206 11554 856
rect 11722 206 11738 856
rect 11906 206 11922 856
rect 12090 206 12198 856
rect 12366 206 12382 856
rect 12550 206 12658 856
rect 12826 206 12842 856
rect 13010 206 13026 856
rect 13194 206 13302 856
rect 13470 206 13486 856
rect 13654 206 13670 856
rect 13838 206 13946 856
rect 14114 206 14130 856
rect 14298 206 14314 856
rect 14482 206 14590 856
rect 14758 206 14774 856
rect 14942 206 15050 856
rect 15218 206 15234 856
rect 15402 206 15418 856
rect 15586 206 15694 856
rect 15862 206 15878 856
rect 16046 206 16062 856
rect 16230 206 16338 856
rect 16506 206 16522 856
rect 16690 206 16706 856
rect 16874 206 16982 856
rect 17150 206 17166 856
rect 17334 206 17442 856
rect 17610 206 17626 856
rect 17794 206 17810 856
rect 17978 206 18086 856
rect 18254 206 18270 856
rect 18438 206 18454 856
rect 18622 206 18730 856
rect 18898 206 18914 856
rect 19082 206 19098 856
rect 19266 206 19374 856
rect 19542 206 19558 856
rect 19726 206 19834 856
rect 20002 206 20018 856
rect 20186 206 20202 856
rect 20370 206 20478 856
rect 20646 206 20662 856
rect 20830 206 20846 856
rect 21014 206 21122 856
rect 21290 206 21306 856
rect 21474 206 21490 856
rect 21658 206 21766 856
rect 21934 206 21950 856
rect 22118 206 22226 856
rect 22394 206 22410 856
rect 22578 206 22594 856
rect 22762 206 22870 856
rect 23038 206 23054 856
rect 23222 206 23238 856
rect 23406 206 23514 856
rect 23682 206 23698 856
rect 23866 206 23882 856
rect 24050 206 24158 856
rect 24326 206 24342 856
rect 24510 206 24618 856
rect 24786 206 24802 856
rect 24970 206 24986 856
rect 25154 206 25262 856
rect 25430 206 25446 856
rect 25614 206 25630 856
rect 25798 206 25906 856
rect 26074 206 26090 856
rect 26258 206 26274 856
rect 26442 206 26550 856
rect 26718 206 26734 856
rect 26902 206 27010 856
rect 27178 206 27194 856
rect 27362 206 27378 856
rect 27546 206 27654 856
rect 27822 206 27838 856
rect 28006 206 28022 856
rect 28190 206 28298 856
rect 28466 206 28482 856
rect 28650 206 28666 856
rect 28834 206 28942 856
rect 29110 206 29126 856
rect 29294 206 29402 856
rect 29570 206 29586 856
rect 29754 206 29770 856
rect 29938 206 30046 856
rect 30214 206 30230 856
rect 30398 206 30414 856
rect 30582 206 30690 856
rect 30858 206 30874 856
rect 31042 206 31058 856
rect 31226 206 31334 856
rect 31502 206 31518 856
rect 31686 206 31794 856
rect 31962 206 31978 856
rect 32146 206 32162 856
rect 32330 206 32438 856
rect 32606 206 32622 856
rect 32790 206 32806 856
rect 32974 206 33082 856
rect 33250 206 33266 856
rect 33434 206 33450 856
rect 33618 206 33726 856
rect 33894 206 33910 856
rect 34078 206 34186 856
rect 34354 206 34370 856
rect 34538 206 34554 856
rect 34722 206 34830 856
rect 34998 206 35014 856
rect 35182 206 35198 856
rect 35366 206 35474 856
rect 35642 206 35658 856
rect 35826 206 35842 856
rect 36010 206 36118 856
rect 36286 206 36302 856
rect 36470 206 36578 856
rect 36746 206 36762 856
rect 36930 206 36946 856
rect 37114 206 37222 856
rect 37390 206 37406 856
rect 37574 206 37590 856
rect 37758 206 37866 856
rect 38034 206 38050 856
rect 38218 206 38234 856
rect 38402 206 38510 856
rect 38678 206 38694 856
rect 38862 206 38970 856
rect 39138 206 39154 856
rect 39322 206 39338 856
rect 39506 206 39614 856
rect 39782 206 39798 856
rect 39966 206 39982 856
rect 40150 206 40258 856
rect 40426 206 40442 856
rect 40610 206 40626 856
rect 40794 206 40902 856
rect 41070 206 41086 856
rect 41254 206 41362 856
rect 41530 206 41546 856
rect 41714 206 41730 856
rect 41898 206 42006 856
rect 42174 206 42190 856
rect 42358 206 42374 856
rect 42542 206 42650 856
rect 42818 206 42834 856
rect 43002 206 43018 856
rect 43186 206 43294 856
rect 43462 206 43478 856
rect 43646 206 43754 856
rect 43922 206 43938 856
rect 44106 206 44122 856
rect 44290 206 44398 856
rect 44566 206 44582 856
rect 44750 206 44766 856
rect 44934 206 45042 856
rect 45210 206 45226 856
rect 45394 206 45410 856
rect 45578 206 45686 856
rect 45854 206 45870 856
rect 46038 206 46054 856
rect 46222 206 46330 856
rect 46498 206 46514 856
rect 46682 206 46790 856
rect 46958 206 46974 856
rect 47142 206 47158 856
rect 47326 206 47434 856
rect 47602 206 47618 856
rect 47786 206 47802 856
rect 47970 206 48078 856
rect 48246 206 48262 856
rect 48430 206 48446 856
rect 48614 206 48722 856
rect 48890 206 48906 856
rect 49074 206 49182 856
rect 49350 206 49366 856
rect 49534 206 49550 856
rect 49718 206 49826 856
rect 49994 206 50010 856
rect 50178 206 50194 856
rect 50362 206 50470 856
rect 50638 206 50654 856
rect 50822 206 50838 856
rect 51006 206 51114 856
rect 51282 206 51298 856
rect 51466 206 51574 856
rect 51742 206 51758 856
rect 51926 206 51942 856
rect 52110 206 52218 856
rect 52386 206 52402 856
rect 52570 206 52586 856
rect 52754 206 52862 856
rect 53030 206 53046 856
rect 53214 206 53230 856
rect 53398 206 53506 856
rect 53674 206 53690 856
rect 53858 206 53966 856
rect 54134 206 54150 856
rect 54318 206 54334 856
rect 54502 206 54610 856
rect 54778 206 54794 856
rect 54962 206 54978 856
rect 55146 206 55254 856
rect 55422 206 55438 856
rect 55606 206 55622 856
rect 55790 206 55898 856
rect 56066 206 56082 856
rect 56250 206 56358 856
rect 56526 206 56542 856
rect 56710 206 56726 856
rect 56894 206 57002 856
rect 57170 206 57186 856
rect 57354 206 57370 856
rect 57538 206 57646 856
rect 57814 206 57830 856
rect 57998 206 58014 856
rect 58182 206 58290 856
rect 58458 206 58474 856
rect 58642 206 58750 856
rect 58918 206 58934 856
rect 59102 206 59118 856
rect 59286 206 59394 856
rect 59562 206 59578 856
rect 59746 206 59762 856
rect 59930 206 60038 856
rect 60206 206 60222 856
rect 60390 206 60406 856
rect 60574 206 60682 856
rect 60850 206 60866 856
rect 61034 206 61142 856
rect 61310 206 61326 856
rect 61494 206 61510 856
rect 61678 206 61786 856
rect 61954 206 61970 856
rect 62138 206 62154 856
rect 62322 206 62430 856
rect 62598 206 62614 856
rect 62782 206 62798 856
rect 62966 206 63074 856
rect 63242 206 63258 856
rect 63426 206 63534 856
rect 63702 206 63718 856
rect 63886 206 63902 856
rect 64070 206 64178 856
rect 64346 206 64362 856
rect 64530 206 64546 856
rect 64714 206 64822 856
rect 64990 206 65006 856
rect 65174 206 65190 856
rect 65358 206 65466 856
rect 65634 206 65650 856
rect 65818 206 65926 856
rect 66094 206 66110 856
rect 66278 206 66294 856
rect 66462 206 66570 856
rect 66738 206 66754 856
rect 66922 206 66938 856
rect 67106 206 67214 856
rect 67382 206 67398 856
rect 67566 206 67582 856
rect 67750 206 67858 856
rect 68026 206 68042 856
rect 68210 206 68318 856
rect 68486 206 68502 856
rect 68670 206 68686 856
rect 68854 206 68962 856
rect 69130 206 69146 856
rect 69314 206 69330 856
rect 69498 206 69606 856
rect 69774 206 69790 856
rect 69958 206 69974 856
rect 70142 206 70250 856
rect 70418 206 70434 856
rect 70602 206 70710 856
rect 70878 206 70894 856
rect 71062 206 71078 856
rect 71246 206 71354 856
rect 71522 206 71538 856
rect 71706 206 71722 856
rect 71890 206 71998 856
rect 72166 206 72182 856
rect 72350 206 72366 856
rect 72534 206 72642 856
rect 72810 206 72826 856
rect 72994 206 73102 856
rect 73270 206 73286 856
rect 73454 206 73470 856
rect 73638 206 73746 856
rect 73914 206 73930 856
rect 74098 206 74114 856
rect 74282 206 74390 856
rect 74558 206 74574 856
rect 74742 206 74758 856
rect 74926 206 75034 856
rect 75202 206 75218 856
rect 75386 206 75494 856
rect 75662 206 75678 856
rect 75846 206 75862 856
rect 76030 206 76138 856
rect 76306 206 76322 856
rect 76490 206 76506 856
rect 76674 206 76782 856
rect 76950 206 76966 856
rect 77134 206 77150 856
rect 77318 206 77426 856
rect 77594 206 77610 856
rect 77778 206 77886 856
rect 78054 206 78070 856
rect 78238 206 78254 856
rect 78422 206 78530 856
rect 78698 206 78714 856
rect 78882 206 78898 856
rect 79066 206 79174 856
rect 79342 206 79358 856
rect 79526 206 79542 856
rect 79710 206 79818 856
rect 79986 206 80002 856
rect 80170 206 80278 856
rect 80446 206 80462 856
rect 80630 206 80646 856
rect 80814 206 80922 856
rect 81090 206 81106 856
rect 81274 206 81290 856
rect 81458 206 81566 856
rect 81734 206 81750 856
rect 81918 206 81934 856
rect 82102 206 82210 856
rect 82378 206 82394 856
rect 82562 206 82670 856
rect 82838 206 82854 856
rect 83022 206 83038 856
rect 83206 206 83314 856
rect 83482 206 83498 856
rect 83666 206 83682 856
rect 83850 206 83958 856
rect 84126 206 84142 856
rect 84310 206 84326 856
rect 84494 206 84602 856
rect 84770 206 84786 856
rect 84954 206 85062 856
rect 85230 206 85246 856
rect 85414 206 85430 856
rect 85598 206 85706 856
rect 85874 206 85890 856
rect 86058 206 86074 856
rect 86242 206 86350 856
rect 86518 206 86534 856
rect 86702 206 86718 856
rect 86886 206 86994 856
rect 87162 206 87178 856
rect 87346 206 87454 856
rect 87622 206 87638 856
rect 87806 206 87822 856
rect 87990 206 88098 856
rect 88266 206 88282 856
rect 88450 206 88466 856
rect 88634 206 88742 856
rect 88910 206 88926 856
rect 89094 206 89110 856
rect 89278 206 89386 856
rect 89554 206 89570 856
rect 89738 206 89754 856
rect 89922 206 90030 856
rect 90198 206 90214 856
rect 90382 206 90490 856
rect 90658 206 90674 856
rect 90842 206 90858 856
rect 91026 206 91134 856
rect 91302 206 91318 856
rect 91486 206 91502 856
rect 91670 206 91778 856
rect 91946 206 91962 856
rect 92130 206 92146 856
rect 92314 206 92422 856
rect 92590 206 92606 856
rect 92774 206 92882 856
rect 93050 206 93066 856
rect 93234 206 93250 856
rect 93418 206 93526 856
rect 93694 206 93710 856
rect 93878 206 93894 856
rect 94062 206 94170 856
rect 94338 206 94354 856
rect 94522 206 94538 856
rect 94706 206 94814 856
rect 94982 206 94998 856
rect 95166 206 95274 856
rect 95442 206 95458 856
rect 95626 206 95642 856
rect 95810 206 95918 856
rect 96086 206 96102 856
rect 96270 206 96286 856
rect 96454 206 96562 856
rect 96730 206 96746 856
rect 96914 206 96930 856
rect 97098 206 97206 856
rect 97374 206 97390 856
rect 97558 206 97666 856
rect 97834 206 97850 856
rect 98018 206 98034 856
rect 98202 206 98310 856
rect 98478 206 98494 856
rect 98662 206 98678 856
rect 98846 206 98954 856
rect 99122 206 99138 856
rect 99306 206 99322 856
rect 99490 206 99598 856
rect 99766 206 99782 856
rect 99950 206 100058 856
rect 100226 206 100242 856
rect 100410 206 100426 856
rect 100594 206 100702 856
rect 100870 206 100886 856
rect 101054 206 101070 856
rect 101238 206 101346 856
rect 101514 206 101530 856
rect 101698 206 101714 856
rect 101882 206 101990 856
rect 102158 206 102174 856
rect 102342 206 102450 856
rect 102618 206 102634 856
rect 102802 206 102818 856
rect 102986 206 103094 856
rect 103262 206 103278 856
rect 103446 206 103462 856
rect 103630 206 103738 856
rect 103906 206 103922 856
rect 104090 206 104106 856
rect 104274 206 104382 856
rect 104550 206 104566 856
rect 104734 206 104842 856
rect 105010 206 105026 856
rect 105194 206 105210 856
rect 105378 206 105486 856
rect 105654 206 105670 856
rect 105838 206 105854 856
rect 106022 206 106130 856
rect 106298 206 106314 856
rect 106482 206 106498 856
rect 106666 206 106774 856
rect 106942 206 106958 856
rect 107126 206 107234 856
rect 107402 206 107418 856
rect 107586 206 107602 856
rect 107770 206 107878 856
rect 108046 206 108062 856
rect 108230 206 108246 856
rect 108414 206 108522 856
rect 108690 206 108706 856
rect 108874 206 108890 856
rect 109058 206 109166 856
rect 109334 206 109350 856
rect 109518 206 109626 856
rect 109794 206 109810 856
rect 109978 206 109994 856
rect 110162 206 110270 856
rect 110438 206 110454 856
rect 110622 206 110638 856
rect 110806 206 110914 856
rect 111082 206 111098 856
rect 111266 206 111282 856
rect 111450 206 111558 856
rect 111726 206 111742 856
rect 111910 206 112018 856
rect 112186 206 112202 856
rect 112370 206 112386 856
rect 112554 206 112662 856
rect 112830 206 112846 856
rect 113014 206 113030 856
rect 113198 206 113306 856
rect 113474 206 113490 856
rect 113658 206 113674 856
rect 113842 206 113950 856
rect 114118 206 114134 856
rect 114302 206 114410 856
rect 114578 206 114594 856
rect 114762 206 114778 856
rect 114946 206 115054 856
rect 115222 206 115238 856
rect 115406 206 115422 856
rect 115590 206 115698 856
rect 115866 206 115882 856
rect 116050 206 116066 856
rect 116234 206 116342 856
rect 116510 206 116526 856
rect 116694 206 116802 856
rect 116970 206 116986 856
rect 117154 206 117170 856
rect 117338 206 117446 856
rect 117614 206 117630 856
rect 117798 206 117814 856
rect 117982 206 118090 856
rect 118258 206 118274 856
rect 118442 206 118458 856
rect 118626 206 118734 856
rect 118902 206 118918 856
rect 119086 206 119194 856
rect 119362 206 119378 856
rect 119546 206 119562 856
rect 119730 206 119838 856
rect 120006 206 120022 856
rect 120190 206 120206 856
rect 120374 206 120482 856
rect 120650 206 120666 856
rect 120834 206 120850 856
rect 121018 206 121126 856
rect 121294 206 121310 856
rect 121478 206 121586 856
rect 121754 206 121770 856
rect 121938 206 121954 856
rect 122122 206 122230 856
rect 122398 206 122414 856
rect 122582 206 122598 856
rect 122766 206 122874 856
rect 123042 206 123058 856
rect 123226 206 123242 856
rect 123410 206 123518 856
rect 123686 206 123702 856
rect 123870 206 123978 856
rect 124146 206 124162 856
rect 124330 206 124346 856
rect 124514 206 124622 856
rect 124790 206 124806 856
rect 124974 206 124990 856
rect 125158 206 125266 856
rect 125434 206 125450 856
rect 125618 206 125634 856
rect 125802 206 125910 856
rect 126078 206 126094 856
rect 126262 206 126370 856
rect 126538 206 126554 856
rect 126722 206 126738 856
rect 126906 206 127014 856
rect 127182 206 127198 856
rect 127366 206 127382 856
rect 127550 206 127658 856
rect 127826 206 127842 856
rect 128010 206 128026 856
rect 128194 206 128302 856
rect 128470 206 128486 856
rect 128654 206 128762 856
rect 128930 206 128946 856
rect 129114 206 129130 856
rect 129298 206 129406 856
rect 129574 206 129590 856
rect 129758 206 129774 856
rect 129942 206 130050 856
rect 130218 206 130234 856
rect 130402 206 130418 856
rect 130586 206 130694 856
rect 130862 206 130878 856
<< obsm3 >>
rect 933 446 129891 130593
<< metal4 >>
rect 4208 2128 4528 130608
rect 19568 2128 19888 130608
rect 34928 2128 35248 130608
rect 50288 2128 50608 130608
rect 65648 2128 65968 130608
rect 81008 2128 81328 130608
rect 96368 2128 96688 130608
rect 111728 2128 112048 130608
rect 127088 2128 127408 130608
<< obsm4 >>
rect 2267 2048 4128 129845
rect 4608 2048 19488 129845
rect 19968 2048 34848 129845
rect 35328 2048 50208 129845
rect 50688 2048 65568 129845
rect 66048 2048 80928 129845
rect 81408 2048 96288 129845
rect 96768 2048 111648 129845
rect 112128 2048 127008 129845
rect 127488 2048 127637 129845
rect 2267 715 127637 2048
<< labels >>
rlabel metal2 s 2686 132408 2742 133208 6 dram_addr0[0]
port 1 nsew signal output
rlabel metal2 s 5814 132408 5870 133208 6 dram_addr0[1]
port 2 nsew signal output
rlabel metal2 s 8850 132408 8906 133208 6 dram_addr0[2]
port 3 nsew signal output
rlabel metal2 s 11978 132408 12034 133208 6 dram_addr0[3]
port 4 nsew signal output
rlabel metal2 s 15106 132408 15162 133208 6 dram_addr0[4]
port 5 nsew signal output
rlabel metal2 s 17406 132408 17462 133208 6 dram_addr0[5]
port 6 nsew signal output
rlabel metal2 s 19706 132408 19762 133208 6 dram_addr0[6]
port 7 nsew signal output
rlabel metal2 s 22098 132408 22154 133208 6 dram_addr0[7]
port 8 nsew signal output
rlabel metal2 s 24398 132408 24454 133208 6 dram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 386 132408 442 133208 6 dram_clk0
port 10 nsew signal output
rlabel metal2 s 1122 132408 1178 133208 6 dram_csb0
port 11 nsew signal output
rlabel metal2 s 3422 132408 3478 133208 6 dram_din0[0]
port 12 nsew signal output
rlabel metal2 s 28262 132408 28318 133208 6 dram_din0[10]
port 13 nsew signal output
rlabel metal2 s 29826 132408 29882 133208 6 dram_din0[11]
port 14 nsew signal output
rlabel metal2 s 31390 132408 31446 133208 6 dram_din0[12]
port 15 nsew signal output
rlabel metal2 s 32954 132408 33010 133208 6 dram_din0[13]
port 16 nsew signal output
rlabel metal2 s 34518 132408 34574 133208 6 dram_din0[14]
port 17 nsew signal output
rlabel metal2 s 35990 132408 36046 133208 6 dram_din0[15]
port 18 nsew signal output
rlabel metal2 s 37554 132408 37610 133208 6 dram_din0[16]
port 19 nsew signal output
rlabel metal2 s 39118 132408 39174 133208 6 dram_din0[17]
port 20 nsew signal output
rlabel metal2 s 40682 132408 40738 133208 6 dram_din0[18]
port 21 nsew signal output
rlabel metal2 s 42246 132408 42302 133208 6 dram_din0[19]
port 22 nsew signal output
rlabel metal2 s 6550 132408 6606 133208 6 dram_din0[1]
port 23 nsew signal output
rlabel metal2 s 43810 132408 43866 133208 6 dram_din0[20]
port 24 nsew signal output
rlabel metal2 s 45374 132408 45430 133208 6 dram_din0[21]
port 25 nsew signal output
rlabel metal2 s 46846 132408 46902 133208 6 dram_din0[22]
port 26 nsew signal output
rlabel metal2 s 48410 132408 48466 133208 6 dram_din0[23]
port 27 nsew signal output
rlabel metal2 s 49974 132408 50030 133208 6 dram_din0[24]
port 28 nsew signal output
rlabel metal2 s 51538 132408 51594 133208 6 dram_din0[25]
port 29 nsew signal output
rlabel metal2 s 53102 132408 53158 133208 6 dram_din0[26]
port 30 nsew signal output
rlabel metal2 s 54666 132408 54722 133208 6 dram_din0[27]
port 31 nsew signal output
rlabel metal2 s 56230 132408 56286 133208 6 dram_din0[28]
port 32 nsew signal output
rlabel metal2 s 57702 132408 57758 133208 6 dram_din0[29]
port 33 nsew signal output
rlabel metal2 s 9678 132408 9734 133208 6 dram_din0[2]
port 34 nsew signal output
rlabel metal2 s 59266 132408 59322 133208 6 dram_din0[30]
port 35 nsew signal output
rlabel metal2 s 60830 132408 60886 133208 6 dram_din0[31]
port 36 nsew signal output
rlabel metal2 s 12714 132408 12770 133208 6 dram_din0[3]
port 37 nsew signal output
rlabel metal2 s 15842 132408 15898 133208 6 dram_din0[4]
port 38 nsew signal output
rlabel metal2 s 18142 132408 18198 133208 6 dram_din0[5]
port 39 nsew signal output
rlabel metal2 s 20534 132408 20590 133208 6 dram_din0[6]
port 40 nsew signal output
rlabel metal2 s 22834 132408 22890 133208 6 dram_din0[7]
port 41 nsew signal output
rlabel metal2 s 25134 132408 25190 133208 6 dram_din0[8]
port 42 nsew signal output
rlabel metal2 s 26698 132408 26754 133208 6 dram_din0[9]
port 43 nsew signal output
rlabel metal2 s 4250 132408 4306 133208 6 dram_dout0[0]
port 44 nsew signal input
rlabel metal2 s 28998 132408 29054 133208 6 dram_dout0[10]
port 45 nsew signal input
rlabel metal2 s 30562 132408 30618 133208 6 dram_dout0[11]
port 46 nsew signal input
rlabel metal2 s 32126 132408 32182 133208 6 dram_dout0[12]
port 47 nsew signal input
rlabel metal2 s 33690 132408 33746 133208 6 dram_dout0[13]
port 48 nsew signal input
rlabel metal2 s 35254 132408 35310 133208 6 dram_dout0[14]
port 49 nsew signal input
rlabel metal2 s 36818 132408 36874 133208 6 dram_dout0[15]
port 50 nsew signal input
rlabel metal2 s 38382 132408 38438 133208 6 dram_dout0[16]
port 51 nsew signal input
rlabel metal2 s 39946 132408 40002 133208 6 dram_dout0[17]
port 52 nsew signal input
rlabel metal2 s 41418 132408 41474 133208 6 dram_dout0[18]
port 53 nsew signal input
rlabel metal2 s 42982 132408 43038 133208 6 dram_dout0[19]
port 54 nsew signal input
rlabel metal2 s 7286 132408 7342 133208 6 dram_dout0[1]
port 55 nsew signal input
rlabel metal2 s 44546 132408 44602 133208 6 dram_dout0[20]
port 56 nsew signal input
rlabel metal2 s 46110 132408 46166 133208 6 dram_dout0[21]
port 57 nsew signal input
rlabel metal2 s 47674 132408 47730 133208 6 dram_dout0[22]
port 58 nsew signal input
rlabel metal2 s 49238 132408 49294 133208 6 dram_dout0[23]
port 59 nsew signal input
rlabel metal2 s 50802 132408 50858 133208 6 dram_dout0[24]
port 60 nsew signal input
rlabel metal2 s 52274 132408 52330 133208 6 dram_dout0[25]
port 61 nsew signal input
rlabel metal2 s 53838 132408 53894 133208 6 dram_dout0[26]
port 62 nsew signal input
rlabel metal2 s 55402 132408 55458 133208 6 dram_dout0[27]
port 63 nsew signal input
rlabel metal2 s 56966 132408 57022 133208 6 dram_dout0[28]
port 64 nsew signal input
rlabel metal2 s 58530 132408 58586 133208 6 dram_dout0[29]
port 65 nsew signal input
rlabel metal2 s 10414 132408 10470 133208 6 dram_dout0[2]
port 66 nsew signal input
rlabel metal2 s 60094 132408 60150 133208 6 dram_dout0[30]
port 67 nsew signal input
rlabel metal2 s 61658 132408 61714 133208 6 dram_dout0[31]
port 68 nsew signal input
rlabel metal2 s 13542 132408 13598 133208 6 dram_dout0[3]
port 69 nsew signal input
rlabel metal2 s 16670 132408 16726 133208 6 dram_dout0[4]
port 70 nsew signal input
rlabel metal2 s 18970 132408 19026 133208 6 dram_dout0[5]
port 71 nsew signal input
rlabel metal2 s 21270 132408 21326 133208 6 dram_dout0[6]
port 72 nsew signal input
rlabel metal2 s 23570 132408 23626 133208 6 dram_dout0[7]
port 73 nsew signal input
rlabel metal2 s 25962 132408 26018 133208 6 dram_dout0[8]
port 74 nsew signal input
rlabel metal2 s 27526 132408 27582 133208 6 dram_dout0[9]
port 75 nsew signal input
rlabel metal2 s 1858 132408 1914 133208 6 dram_web0
port 76 nsew signal output
rlabel metal2 s 4986 132408 5042 133208 6 dram_wmask0[0]
port 77 nsew signal output
rlabel metal2 s 8114 132408 8170 133208 6 dram_wmask0[1]
port 78 nsew signal output
rlabel metal2 s 11242 132408 11298 133208 6 dram_wmask0[2]
port 79 nsew signal output
rlabel metal2 s 14278 132408 14334 133208 6 dram_wmask0[3]
port 80 nsew signal output
rlabel metal2 s 64694 132408 64750 133208 6 gpio_in[0]
port 81 nsew signal input
rlabel metal2 s 87970 132408 88026 133208 6 gpio_in[10]
port 82 nsew signal input
rlabel metal2 s 90362 132408 90418 133208 6 gpio_in[11]
port 83 nsew signal input
rlabel metal2 s 92662 132408 92718 133208 6 gpio_in[12]
port 84 nsew signal input
rlabel metal2 s 94962 132408 95018 133208 6 gpio_in[13]
port 85 nsew signal input
rlabel metal2 s 97262 132408 97318 133208 6 gpio_in[14]
port 86 nsew signal input
rlabel metal2 s 99654 132408 99710 133208 6 gpio_in[15]
port 87 nsew signal input
rlabel metal2 s 101954 132408 102010 133208 6 gpio_in[16]
port 88 nsew signal input
rlabel metal2 s 104254 132408 104310 133208 6 gpio_in[17]
port 89 nsew signal input
rlabel metal2 s 106646 132408 106702 133208 6 gpio_in[18]
port 90 nsew signal input
rlabel metal2 s 108946 132408 109002 133208 6 gpio_in[19]
port 91 nsew signal input
rlabel metal2 s 67086 132408 67142 133208 6 gpio_in[1]
port 92 nsew signal input
rlabel metal2 s 111246 132408 111302 133208 6 gpio_in[20]
port 93 nsew signal input
rlabel metal2 s 113638 132408 113694 133208 6 gpio_in[21]
port 94 nsew signal input
rlabel metal2 s 115938 132408 115994 133208 6 gpio_in[22]
port 95 nsew signal input
rlabel metal2 s 118238 132408 118294 133208 6 gpio_in[23]
port 96 nsew signal input
rlabel metal2 s 69386 132408 69442 133208 6 gpio_in[2]
port 97 nsew signal input
rlabel metal2 s 71686 132408 71742 133208 6 gpio_in[3]
port 98 nsew signal input
rlabel metal2 s 74078 132408 74134 133208 6 gpio_in[4]
port 99 nsew signal input
rlabel metal2 s 76378 132408 76434 133208 6 gpio_in[5]
port 100 nsew signal input
rlabel metal2 s 78678 132408 78734 133208 6 gpio_in[6]
port 101 nsew signal input
rlabel metal2 s 80978 132408 81034 133208 6 gpio_in[7]
port 102 nsew signal input
rlabel metal2 s 83370 132408 83426 133208 6 gpio_in[8]
port 103 nsew signal input
rlabel metal2 s 85670 132408 85726 133208 6 gpio_in[9]
port 104 nsew signal input
rlabel metal2 s 65522 132408 65578 133208 6 gpio_oeb[0]
port 105 nsew signal output
rlabel metal2 s 88798 132408 88854 133208 6 gpio_oeb[10]
port 106 nsew signal output
rlabel metal2 s 91098 132408 91154 133208 6 gpio_oeb[11]
port 107 nsew signal output
rlabel metal2 s 93398 132408 93454 133208 6 gpio_oeb[12]
port 108 nsew signal output
rlabel metal2 s 95790 132408 95846 133208 6 gpio_oeb[13]
port 109 nsew signal output
rlabel metal2 s 98090 132408 98146 133208 6 gpio_oeb[14]
port 110 nsew signal output
rlabel metal2 s 100390 132408 100446 133208 6 gpio_oeb[15]
port 111 nsew signal output
rlabel metal2 s 102782 132408 102838 133208 6 gpio_oeb[16]
port 112 nsew signal output
rlabel metal2 s 105082 132408 105138 133208 6 gpio_oeb[17]
port 113 nsew signal output
rlabel metal2 s 107382 132408 107438 133208 6 gpio_oeb[18]
port 114 nsew signal output
rlabel metal2 s 109682 132408 109738 133208 6 gpio_oeb[19]
port 115 nsew signal output
rlabel metal2 s 67822 132408 67878 133208 6 gpio_oeb[1]
port 116 nsew signal output
rlabel metal2 s 112074 132408 112130 133208 6 gpio_oeb[20]
port 117 nsew signal output
rlabel metal2 s 114374 132408 114430 133208 6 gpio_oeb[21]
port 118 nsew signal output
rlabel metal2 s 116674 132408 116730 133208 6 gpio_oeb[22]
port 119 nsew signal output
rlabel metal2 s 119066 132408 119122 133208 6 gpio_oeb[23]
port 120 nsew signal output
rlabel metal2 s 120538 132408 120594 133208 6 gpio_oeb[24]
port 121 nsew signal output
rlabel metal2 s 121366 132408 121422 133208 6 gpio_oeb[25]
port 122 nsew signal output
rlabel metal2 s 122102 132408 122158 133208 6 gpio_oeb[26]
port 123 nsew signal output
rlabel metal2 s 122930 132408 122986 133208 6 gpio_oeb[27]
port 124 nsew signal output
rlabel metal2 s 123666 132408 123722 133208 6 gpio_oeb[28]
port 125 nsew signal output
rlabel metal2 s 124494 132408 124550 133208 6 gpio_oeb[29]
port 126 nsew signal output
rlabel metal2 s 70122 132408 70178 133208 6 gpio_oeb[2]
port 127 nsew signal output
rlabel metal2 s 125230 132408 125286 133208 6 gpio_oeb[30]
port 128 nsew signal output
rlabel metal2 s 125966 132408 126022 133208 6 gpio_oeb[31]
port 129 nsew signal output
rlabel metal2 s 126794 132408 126850 133208 6 gpio_oeb[32]
port 130 nsew signal output
rlabel metal2 s 127530 132408 127586 133208 6 gpio_oeb[33]
port 131 nsew signal output
rlabel metal2 s 128358 132408 128414 133208 6 gpio_oeb[34]
port 132 nsew signal output
rlabel metal2 s 129094 132408 129150 133208 6 gpio_oeb[35]
port 133 nsew signal output
rlabel metal2 s 129922 132408 129978 133208 6 gpio_oeb[36]
port 134 nsew signal output
rlabel metal2 s 130658 132408 130714 133208 6 gpio_oeb[37]
port 135 nsew signal output
rlabel metal2 s 72514 132408 72570 133208 6 gpio_oeb[3]
port 136 nsew signal output
rlabel metal2 s 74814 132408 74870 133208 6 gpio_oeb[4]
port 137 nsew signal output
rlabel metal2 s 77114 132408 77170 133208 6 gpio_oeb[5]
port 138 nsew signal output
rlabel metal2 s 79506 132408 79562 133208 6 gpio_oeb[6]
port 139 nsew signal output
rlabel metal2 s 81806 132408 81862 133208 6 gpio_oeb[7]
port 140 nsew signal output
rlabel metal2 s 84106 132408 84162 133208 6 gpio_oeb[8]
port 141 nsew signal output
rlabel metal2 s 86406 132408 86462 133208 6 gpio_oeb[9]
port 142 nsew signal output
rlabel metal2 s 66258 132408 66314 133208 6 gpio_out[0]
port 143 nsew signal output
rlabel metal2 s 89534 132408 89590 133208 6 gpio_out[10]
port 144 nsew signal output
rlabel metal2 s 91834 132408 91890 133208 6 gpio_out[11]
port 145 nsew signal output
rlabel metal2 s 94226 132408 94282 133208 6 gpio_out[12]
port 146 nsew signal output
rlabel metal2 s 96526 132408 96582 133208 6 gpio_out[13]
port 147 nsew signal output
rlabel metal2 s 98826 132408 98882 133208 6 gpio_out[14]
port 148 nsew signal output
rlabel metal2 s 101218 132408 101274 133208 6 gpio_out[15]
port 149 nsew signal output
rlabel metal2 s 103518 132408 103574 133208 6 gpio_out[16]
port 150 nsew signal output
rlabel metal2 s 105818 132408 105874 133208 6 gpio_out[17]
port 151 nsew signal output
rlabel metal2 s 108210 132408 108266 133208 6 gpio_out[18]
port 152 nsew signal output
rlabel metal2 s 110510 132408 110566 133208 6 gpio_out[19]
port 153 nsew signal output
rlabel metal2 s 68650 132408 68706 133208 6 gpio_out[1]
port 154 nsew signal output
rlabel metal2 s 112810 132408 112866 133208 6 gpio_out[20]
port 155 nsew signal output
rlabel metal2 s 115110 132408 115166 133208 6 gpio_out[21]
port 156 nsew signal output
rlabel metal2 s 117502 132408 117558 133208 6 gpio_out[22]
port 157 nsew signal output
rlabel metal2 s 119802 132408 119858 133208 6 gpio_out[23]
port 158 nsew signal output
rlabel metal2 s 70950 132408 71006 133208 6 gpio_out[2]
port 159 nsew signal output
rlabel metal2 s 73250 132408 73306 133208 6 gpio_out[3]
port 160 nsew signal output
rlabel metal2 s 75550 132408 75606 133208 6 gpio_out[4]
port 161 nsew signal output
rlabel metal2 s 77942 132408 77998 133208 6 gpio_out[5]
port 162 nsew signal output
rlabel metal2 s 80242 132408 80298 133208 6 gpio_out[6]
port 163 nsew signal output
rlabel metal2 s 82542 132408 82598 133208 6 gpio_out[7]
port 164 nsew signal output
rlabel metal2 s 84934 132408 84990 133208 6 gpio_out[8]
port 165 nsew signal output
rlabel metal2 s 87234 132408 87290 133208 6 gpio_out[9]
port 166 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 iram_addr0[0]
port 167 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 iram_addr0[1]
port 168 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 iram_addr0[2]
port 169 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 iram_addr0[3]
port 170 nsew signal output
rlabel metal2 s 111798 0 111854 800 6 iram_addr0[4]
port 171 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 iram_addr0[5]
port 172 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 iram_addr0[6]
port 173 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 iram_addr0[7]
port 174 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 iram_addr0[8]
port 175 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 iram_clk0
port 176 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 iram_csb0_A
port 177 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 iram_csb0_B
port 178 nsew signal output
rlabel metal2 s 107658 0 107714 800 6 iram_din0[0]
port 179 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 iram_din0[10]
port 180 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 iram_din0[11]
port 181 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 iram_din0[12]
port 182 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 iram_din0[13]
port 183 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 iram_din0[14]
port 184 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 iram_din0[15]
port 185 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 iram_din0[16]
port 186 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 iram_din0[17]
port 187 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 iram_din0[18]
port 188 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 iram_din0[19]
port 189 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 iram_din0[1]
port 190 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 iram_din0[20]
port 191 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 iram_din0[21]
port 192 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 iram_din0[22]
port 193 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 iram_din0[23]
port 194 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 iram_din0[24]
port 195 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 iram_din0[25]
port 196 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 iram_din0[26]
port 197 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 iram_din0[27]
port 198 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 iram_din0[28]
port 199 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 iram_din0[29]
port 200 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 iram_din0[2]
port 201 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 iram_din0[30]
port 202 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 iram_din0[31]
port 203 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 iram_din0[3]
port 204 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 iram_din0[4]
port 205 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 iram_din0[5]
port 206 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 iram_din0[6]
port 207 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 iram_din0[7]
port 208 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 iram_din0[8]
port 209 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 iram_din0[9]
port 210 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 iram_dout0_A[0]
port 211 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 iram_dout0_A[10]
port 212 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 iram_dout0_A[11]
port 213 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 iram_dout0_A[12]
port 214 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 iram_dout0_A[13]
port 215 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 iram_dout0_A[14]
port 216 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 iram_dout0_A[15]
port 217 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 iram_dout0_A[16]
port 218 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 iram_dout0_A[17]
port 219 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 iram_dout0_A[18]
port 220 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 iram_dout0_A[19]
port 221 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 iram_dout0_A[1]
port 222 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 iram_dout0_A[20]
port 223 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 iram_dout0_A[21]
port 224 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 iram_dout0_A[22]
port 225 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 iram_dout0_A[23]
port 226 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 iram_dout0_A[24]
port 227 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 iram_dout0_A[25]
port 228 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 iram_dout0_A[26]
port 229 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 iram_dout0_A[27]
port 230 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 iram_dout0_A[28]
port 231 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 iram_dout0_A[29]
port 232 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 iram_dout0_A[2]
port 233 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 iram_dout0_A[30]
port 234 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 iram_dout0_A[31]
port 235 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 iram_dout0_A[3]
port 236 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 iram_dout0_A[4]
port 237 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 iram_dout0_A[5]
port 238 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 iram_dout0_A[6]
port 239 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 iram_dout0_A[7]
port 240 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 iram_dout0_A[8]
port 241 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 iram_dout0_A[9]
port 242 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 iram_dout0_B[0]
port 243 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 iram_dout0_B[10]
port 244 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 iram_dout0_B[11]
port 245 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 iram_dout0_B[12]
port 246 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 iram_dout0_B[13]
port 247 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 iram_dout0_B[14]
port 248 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 iram_dout0_B[15]
port 249 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 iram_dout0_B[16]
port 250 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 iram_dout0_B[17]
port 251 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 iram_dout0_B[18]
port 252 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 iram_dout0_B[19]
port 253 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 iram_dout0_B[1]
port 254 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 iram_dout0_B[20]
port 255 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 iram_dout0_B[21]
port 256 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 iram_dout0_B[22]
port 257 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 iram_dout0_B[23]
port 258 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 iram_dout0_B[24]
port 259 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 iram_dout0_B[25]
port 260 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 iram_dout0_B[26]
port 261 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 iram_dout0_B[27]
port 262 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 iram_dout0_B[28]
port 263 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 iram_dout0_B[29]
port 264 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 iram_dout0_B[2]
port 265 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 iram_dout0_B[30]
port 266 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 iram_dout0_B[31]
port 267 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 iram_dout0_B[3]
port 268 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 iram_dout0_B[4]
port 269 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 iram_dout0_B[5]
port 270 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 iram_dout0_B[6]
port 271 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 iram_dout0_B[7]
port 272 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 iram_dout0_B[8]
port 273 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 iram_dout0_B[9]
port 274 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 iram_web0
port 275 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 iram_wmask0[0]
port 276 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 iram_wmask0[1]
port 277 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 iram_wmask0[2]
port 278 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 iram_wmask0[3]
port 279 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 la_data_in[0]
port 280 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[100]
port 281 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[101]
port 282 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_data_in[102]
port 283 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[103]
port 284 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[104]
port 285 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[105]
port 286 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[106]
port 287 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[107]
port 288 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[108]
port 289 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[109]
port 290 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_data_in[10]
port 291 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[110]
port 292 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[111]
port 293 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[112]
port 294 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[113]
port 295 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[114]
port 296 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_data_in[115]
port 297 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[116]
port 298 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[117]
port 299 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[118]
port 300 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[119]
port 301 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[11]
port 302 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[120]
port 303 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[121]
port 304 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[122]
port 305 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_data_in[123]
port 306 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[124]
port 307 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[125]
port 308 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[126]
port 309 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_data_in[127]
port 310 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[12]
port 311 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[13]
port 312 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_data_in[14]
port 313 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[15]
port 314 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in[16]
port 315 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[17]
port 316 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in[18]
port 317 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_data_in[19]
port 318 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_data_in[1]
port 319 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_data_in[20]
port 320 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[21]
port 321 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[22]
port 322 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[23]
port 323 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_in[24]
port 324 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_in[25]
port 325 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[26]
port 326 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[27]
port 327 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[28]
port 328 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_data_in[29]
port 329 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_data_in[2]
port 330 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_data_in[30]
port 331 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[31]
port 332 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_data_in[32]
port 333 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[33]
port 334 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[34]
port 335 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[35]
port 336 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[36]
port 337 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[37]
port 338 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[38]
port 339 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[39]
port 340 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_data_in[3]
port 341 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[40]
port 342 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_data_in[41]
port 343 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[42]
port 344 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[43]
port 345 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[44]
port 346 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[45]
port 347 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[46]
port 348 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[47]
port 349 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[48]
port 350 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[49]
port 351 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[4]
port 352 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[50]
port 353 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_data_in[51]
port 354 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[52]
port 355 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[53]
port 356 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[54]
port 357 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[55]
port 358 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[56]
port 359 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[57]
port 360 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[58]
port 361 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[59]
port 362 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_data_in[5]
port 363 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[60]
port 364 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[61]
port 365 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[62]
port 366 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[63]
port 367 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[64]
port 368 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[65]
port 369 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[66]
port 370 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[67]
port 371 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[68]
port 372 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[69]
port 373 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[6]
port 374 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[70]
port 375 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_data_in[71]
port 376 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[72]
port 377 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_data_in[73]
port 378 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[74]
port 379 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[75]
port 380 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[76]
port 381 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[77]
port 382 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[78]
port 383 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[79]
port 384 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[7]
port 385 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[80]
port 386 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[81]
port 387 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_data_in[82]
port 388 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[83]
port 389 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[84]
port 390 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[85]
port 391 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[86]
port 392 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_data_in[87]
port 393 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[88]
port 394 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[89]
port 395 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[8]
port 396 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[90]
port 397 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[91]
port 398 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[92]
port 399 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[93]
port 400 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[94]
port 401 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[95]
port 402 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[96]
port 403 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[97]
port 404 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[98]
port 405 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[99]
port 406 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[9]
port 407 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_data_out[0]
port 408 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[100]
port 409 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[101]
port 410 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[102]
port 411 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[103]
port 412 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[104]
port 413 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[105]
port 414 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[106]
port 415 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[107]
port 416 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[108]
port 417 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[109]
port 418 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 la_data_out[10]
port 419 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[110]
port 420 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[111]
port 421 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[112]
port 422 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[113]
port 423 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[114]
port 424 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[115]
port 425 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[116]
port 426 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 la_data_out[117]
port 427 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[118]
port 428 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[119]
port 429 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 la_data_out[11]
port 430 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[120]
port 431 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[121]
port 432 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[122]
port 433 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[123]
port 434 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[124]
port 435 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[125]
port 436 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[126]
port 437 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[127]
port 438 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 la_data_out[12]
port 439 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 la_data_out[13]
port 440 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 la_data_out[14]
port 441 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 la_data_out[15]
port 442 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_data_out[16]
port 443 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 la_data_out[17]
port 444 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_data_out[18]
port 445 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 la_data_out[19]
port 446 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 la_data_out[1]
port 447 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[20]
port 448 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 la_data_out[21]
port 449 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[22]
port 450 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[23]
port 451 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 la_data_out[24]
port 452 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[25]
port 453 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 la_data_out[26]
port 454 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[27]
port 455 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[28]
port 456 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 la_data_out[29]
port 457 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 la_data_out[2]
port 458 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[30]
port 459 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[31]
port 460 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_data_out[32]
port 461 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[33]
port 462 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[34]
port 463 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[35]
port 464 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[36]
port 465 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[37]
port 466 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[38]
port 467 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[39]
port 468 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[3]
port 469 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[40]
port 470 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[41]
port 471 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[42]
port 472 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_out[43]
port 473 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[44]
port 474 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[45]
port 475 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[46]
port 476 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[47]
port 477 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[48]
port 478 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[49]
port 479 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 la_data_out[4]
port 480 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[50]
port 481 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[51]
port 482 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[52]
port 483 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[53]
port 484 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[54]
port 485 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[55]
port 486 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[56]
port 487 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[57]
port 488 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[58]
port 489 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[59]
port 490 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 la_data_out[5]
port 491 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[60]
port 492 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[61]
port 493 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[62]
port 494 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 la_data_out[63]
port 495 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[64]
port 496 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[65]
port 497 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[66]
port 498 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[67]
port 499 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[68]
port 500 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[69]
port 501 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 la_data_out[6]
port 502 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[70]
port 503 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 la_data_out[71]
port 504 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[72]
port 505 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 la_data_out[73]
port 506 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[74]
port 507 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[75]
port 508 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[76]
port 509 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[77]
port 510 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[78]
port 511 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[79]
port 512 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 la_data_out[7]
port 513 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[80]
port 514 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[81]
port 515 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[82]
port 516 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[83]
port 517 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[84]
port 518 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[85]
port 519 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[86]
port 520 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[87]
port 521 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[88]
port 522 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[89]
port 523 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 la_data_out[8]
port 524 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[90]
port 525 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[91]
port 526 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[92]
port 527 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[93]
port 528 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[94]
port 529 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[95]
port 530 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[96]
port 531 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 la_data_out[97]
port 532 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[98]
port 533 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[99]
port 534 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[9]
port 535 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_oenb[0]
port 536 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[100]
port 537 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_oenb[101]
port 538 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[102]
port 539 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[103]
port 540 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[104]
port 541 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[105]
port 542 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[106]
port 543 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[107]
port 544 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[108]
port 545 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[109]
port 546 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_oenb[10]
port 547 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[110]
port 548 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[111]
port 549 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[112]
port 550 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[113]
port 551 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[114]
port 552 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[115]
port 553 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[116]
port 554 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[117]
port 555 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_oenb[118]
port 556 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[119]
port 557 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_oenb[11]
port 558 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[120]
port 559 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[121]
port 560 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_oenb[122]
port 561 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[123]
port 562 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[124]
port 563 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oenb[125]
port 564 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_oenb[126]
port 565 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_oenb[127]
port 566 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_oenb[12]
port 567 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_oenb[13]
port 568 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_oenb[14]
port 569 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[15]
port 570 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_oenb[16]
port 571 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_oenb[17]
port 572 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[18]
port 573 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[19]
port 574 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_oenb[1]
port 575 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_oenb[20]
port 576 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[21]
port 577 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_oenb[22]
port 578 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_oenb[23]
port 579 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_oenb[24]
port 580 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[25]
port 581 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oenb[26]
port 582 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[27]
port 583 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_oenb[28]
port 584 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[29]
port 585 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_oenb[2]
port 586 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[30]
port 587 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[31]
port 588 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[32]
port 589 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[33]
port 590 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[34]
port 591 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[35]
port 592 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[36]
port 593 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[37]
port 594 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[38]
port 595 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_oenb[39]
port 596 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[3]
port 597 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[40]
port 598 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[41]
port 599 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[42]
port 600 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[43]
port 601 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[44]
port 602 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[45]
port 603 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[46]
port 604 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[47]
port 605 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[48]
port 606 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_oenb[49]
port 607 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_oenb[4]
port 608 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[50]
port 609 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[51]
port 610 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[52]
port 611 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[53]
port 612 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[54]
port 613 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[55]
port 614 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_oenb[56]
port 615 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_oenb[57]
port 616 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[58]
port 617 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_oenb[59]
port 618 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_oenb[5]
port 619 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[60]
port 620 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[61]
port 621 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[62]
port 622 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[63]
port 623 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[64]
port 624 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[65]
port 625 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[66]
port 626 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[67]
port 627 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_oenb[68]
port 628 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[69]
port 629 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_oenb[6]
port 630 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[70]
port 631 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oenb[71]
port 632 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_oenb[72]
port 633 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[73]
port 634 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_oenb[74]
port 635 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[75]
port 636 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_oenb[76]
port 637 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[77]
port 638 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[78]
port 639 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[79]
port 640 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[7]
port 641 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_oenb[80]
port 642 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[81]
port 643 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[82]
port 644 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[83]
port 645 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[84]
port 646 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[85]
port 647 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[86]
port 648 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[87]
port 649 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[88]
port 650 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[89]
port 651 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[8]
port 652 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_oenb[90]
port 653 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_oenb[91]
port 654 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_oenb[92]
port 655 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[93]
port 656 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[94]
port 657 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oenb[95]
port 658 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_oenb[96]
port 659 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[97]
port 660 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[98]
port 661 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[99]
port 662 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_oenb[9]
port 663 nsew signal input
rlabel metal2 s 62394 132408 62450 133208 6 user_irq[0]
port 664 nsew signal output
rlabel metal2 s 63130 132408 63186 133208 6 user_irq[1]
port 665 nsew signal output
rlabel metal2 s 63958 132408 64014 133208 6 user_irq[2]
port 666 nsew signal output
rlabel metal4 s 4208 2128 4528 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 669 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 670 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 671 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[0]
port 672 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[10]
port 673 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[11]
port 674 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[12]
port 675 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_adr_i[13]
port 676 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[14]
port 677 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[15]
port 678 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[16]
port 679 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[17]
port 680 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[18]
port 681 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[19]
port 682 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[1]
port 683 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_adr_i[20]
port 684 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[21]
port 685 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[22]
port 686 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[23]
port 687 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[24]
port 688 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[25]
port 689 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[26]
port 690 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[27]
port 691 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[28]
port 692 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[29]
port 693 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_adr_i[2]
port 694 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[30]
port 695 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[31]
port 696 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[3]
port 697 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[4]
port 698 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[5]
port 699 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[6]
port 700 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[7]
port 701 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[8]
port 702 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[9]
port 703 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 704 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_i[0]
port 705 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[10]
port 706 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[11]
port 707 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[12]
port 708 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[13]
port 709 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[14]
port 710 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[15]
port 711 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[16]
port 712 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_i[17]
port 713 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_i[18]
port 714 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[19]
port 715 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_i[1]
port 716 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_i[20]
port 717 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[21]
port 718 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[22]
port 719 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[23]
port 720 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[24]
port 721 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[25]
port 722 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[26]
port 723 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_i[27]
port 724 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_i[28]
port 725 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[29]
port 726 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[2]
port 727 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[30]
port 728 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[31]
port 729 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[3]
port 730 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_i[4]
port 731 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[5]
port 732 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[6]
port 733 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[7]
port 734 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[8]
port 735 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[9]
port 736 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_o[0]
port 737 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[10]
port 738 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[11]
port 739 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[12]
port 740 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[13]
port 741 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[14]
port 742 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[15]
port 743 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[16]
port 744 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[17]
port 745 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[18]
port 746 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_o[19]
port 747 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[1]
port 748 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_o[20]
port 749 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[21]
port 750 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[22]
port 751 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[23]
port 752 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[24]
port 753 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[25]
port 754 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[26]
port 755 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[27]
port 756 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[28]
port 757 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[29]
port 758 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_o[2]
port 759 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[30]
port 760 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[31]
port 761 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[3]
port 762 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_o[4]
port 763 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[5]
port 764 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[6]
port 765 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[7]
port 766 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[8]
port 767 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[9]
port 768 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 wbs_sel_i[0]
port 769 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_sel_i[1]
port 770 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[2]
port 771 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_sel_i[3]
port 772 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_stb_i
port 773 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 774 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 131064 133208
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 43434258
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc/openlane/rvj1_caravel_soc/runs/rvj1_caravel_soc/results/signoff/rvj1_caravel_soc.magic.gds
string GDS_START 1257002
<< end >>

