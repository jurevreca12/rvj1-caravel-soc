VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wbuart_wrap
  CLASS BLOCK ;
  FOREIGN wbuart_wrap ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.100 BY 360.820 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 251.640 350.100 252.240 ;
    END
  END clk_i
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 356.820 325.590 360.820 ;
    END
  END rst_i
  PIN uart_rx_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 356.820 209.670 360.820 ;
    END
  END uart_rx_i
  PIN uart_tx_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END uart_tx_o
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 348.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 348.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 348.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 348.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 348.400 ;
    END
  END vssd1
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 356.820 196.790 360.820 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 6.840 350.100 7.440 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 306.040 350.100 306.640 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 356.820 145.270 360.820 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 356.820 171.030 360.820 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 129.240 350.100 129.840 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 356.820 248.310 360.820 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 356.820 299.830 360.820 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 346.840 350.100 347.440 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 88.440 350.100 89.040 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 74.840 350.100 75.440 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 61.240 350.100 61.840 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 356.820 183.910 360.820 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 356.820 222.550 360.820 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 278.840 350.100 279.440 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 319.640 350.100 320.240 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 356.820 348.130 360.820 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 356.820 106.630 360.820 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 156.440 350.100 157.040 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 356.820 119.510 360.820 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 292.440 350.100 293.040 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 356.820 132.390 360.820 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 20.440 350.100 21.040 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 197.240 350.100 197.840 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 356.820 80.870 360.820 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 34.040 350.100 34.640 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 333.240 350.100 333.840 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 356.820 286.950 360.820 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 102.040 350.100 102.640 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 356.820 93.750 360.820 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 183.640 350.100 184.240 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 115.640 350.100 116.240 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 142.840 350.100 143.440 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 238.040 350.100 238.640 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 265.240 350.100 265.840 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 356.820 29.350 360.820 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 356.820 42.230 360.820 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 356.820 55.110 360.820 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 356.820 158.150 360.820 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 356.820 312.710 360.820 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 356.820 235.430 360.820 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 356.820 338.470 360.820 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 47.640 350.100 48.240 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 356.820 3.590 360.820 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 210.840 350.100 211.440 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 224.440 350.100 225.040 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 356.820 274.070 360.820 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 356.820 261.190 360.820 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 356.820 16.470 360.820 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 356.820 67.990 360.820 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.100 170.040 350.100 170.640 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.540 348.245 ;
      LAYER met1 ;
        RECT 0.070 9.900 348.150 348.400 ;
      LAYER met2 ;
        RECT 0.100 356.540 3.030 357.410 ;
        RECT 3.870 356.540 15.910 357.410 ;
        RECT 16.750 356.540 28.790 357.410 ;
        RECT 29.630 356.540 41.670 357.410 ;
        RECT 42.510 356.540 54.550 357.410 ;
        RECT 55.390 356.540 67.430 357.410 ;
        RECT 68.270 356.540 80.310 357.410 ;
        RECT 81.150 356.540 93.190 357.410 ;
        RECT 94.030 356.540 106.070 357.410 ;
        RECT 106.910 356.540 118.950 357.410 ;
        RECT 119.790 356.540 131.830 357.410 ;
        RECT 132.670 356.540 144.710 357.410 ;
        RECT 145.550 356.540 157.590 357.410 ;
        RECT 158.430 356.540 170.470 357.410 ;
        RECT 171.310 356.540 183.350 357.410 ;
        RECT 184.190 356.540 196.230 357.410 ;
        RECT 197.070 356.540 209.110 357.410 ;
        RECT 209.950 356.540 221.990 357.410 ;
        RECT 222.830 356.540 234.870 357.410 ;
        RECT 235.710 356.540 247.750 357.410 ;
        RECT 248.590 356.540 260.630 357.410 ;
        RECT 261.470 356.540 273.510 357.410 ;
        RECT 274.350 356.540 286.390 357.410 ;
        RECT 287.230 356.540 299.270 357.410 ;
        RECT 300.110 356.540 312.150 357.410 ;
        RECT 312.990 356.540 325.030 357.410 ;
        RECT 325.870 356.540 337.910 357.410 ;
        RECT 338.750 356.540 347.570 357.410 ;
        RECT 0.100 4.280 348.120 356.540 ;
        RECT 0.650 3.670 9.470 4.280 ;
        RECT 10.310 3.670 22.350 4.280 ;
        RECT 23.190 3.670 35.230 4.280 ;
        RECT 36.070 3.670 48.110 4.280 ;
        RECT 48.950 3.670 60.990 4.280 ;
        RECT 61.830 3.670 73.870 4.280 ;
        RECT 74.710 3.670 86.750 4.280 ;
        RECT 87.590 3.670 99.630 4.280 ;
        RECT 100.470 3.670 112.510 4.280 ;
        RECT 113.350 3.670 125.390 4.280 ;
        RECT 126.230 3.670 138.270 4.280 ;
        RECT 139.110 3.670 151.150 4.280 ;
        RECT 151.990 3.670 164.030 4.280 ;
        RECT 164.870 3.670 176.910 4.280 ;
        RECT 177.750 3.670 189.790 4.280 ;
        RECT 190.630 3.670 202.670 4.280 ;
        RECT 203.510 3.670 215.550 4.280 ;
        RECT 216.390 3.670 228.430 4.280 ;
        RECT 229.270 3.670 241.310 4.280 ;
        RECT 242.150 3.670 254.190 4.280 ;
        RECT 255.030 3.670 267.070 4.280 ;
        RECT 267.910 3.670 279.950 4.280 ;
        RECT 280.790 3.670 292.830 4.280 ;
        RECT 293.670 3.670 305.710 4.280 ;
        RECT 306.550 3.670 318.590 4.280 ;
        RECT 319.430 3.670 331.470 4.280 ;
        RECT 332.310 3.670 344.350 4.280 ;
        RECT 345.190 3.670 348.120 4.280 ;
      LAYER met3 ;
        RECT 4.400 349.840 346.100 350.705 ;
        RECT 4.000 347.840 346.100 349.840 ;
        RECT 4.000 346.440 345.700 347.840 ;
        RECT 4.000 337.640 346.100 346.440 ;
        RECT 4.400 336.240 346.100 337.640 ;
        RECT 4.000 334.240 346.100 336.240 ;
        RECT 4.000 332.840 345.700 334.240 ;
        RECT 4.000 324.040 346.100 332.840 ;
        RECT 4.400 322.640 346.100 324.040 ;
        RECT 4.000 320.640 346.100 322.640 ;
        RECT 4.000 319.240 345.700 320.640 ;
        RECT 4.000 310.440 346.100 319.240 ;
        RECT 4.400 309.040 346.100 310.440 ;
        RECT 4.000 307.040 346.100 309.040 ;
        RECT 4.000 305.640 345.700 307.040 ;
        RECT 4.000 296.840 346.100 305.640 ;
        RECT 4.400 295.440 346.100 296.840 ;
        RECT 4.000 293.440 346.100 295.440 ;
        RECT 4.000 292.040 345.700 293.440 ;
        RECT 4.000 283.240 346.100 292.040 ;
        RECT 4.400 281.840 346.100 283.240 ;
        RECT 4.000 279.840 346.100 281.840 ;
        RECT 4.000 278.440 345.700 279.840 ;
        RECT 4.000 269.640 346.100 278.440 ;
        RECT 4.400 268.240 346.100 269.640 ;
        RECT 4.000 266.240 346.100 268.240 ;
        RECT 4.000 264.840 345.700 266.240 ;
        RECT 4.000 256.040 346.100 264.840 ;
        RECT 4.400 254.640 346.100 256.040 ;
        RECT 4.000 252.640 346.100 254.640 ;
        RECT 4.000 251.240 345.700 252.640 ;
        RECT 4.000 242.440 346.100 251.240 ;
        RECT 4.400 241.040 346.100 242.440 ;
        RECT 4.000 239.040 346.100 241.040 ;
        RECT 4.000 237.640 345.700 239.040 ;
        RECT 4.000 228.840 346.100 237.640 ;
        RECT 4.400 227.440 346.100 228.840 ;
        RECT 4.000 225.440 346.100 227.440 ;
        RECT 4.000 224.040 345.700 225.440 ;
        RECT 4.000 215.240 346.100 224.040 ;
        RECT 4.400 213.840 346.100 215.240 ;
        RECT 4.000 211.840 346.100 213.840 ;
        RECT 4.000 210.440 345.700 211.840 ;
        RECT 4.000 201.640 346.100 210.440 ;
        RECT 4.400 200.240 346.100 201.640 ;
        RECT 4.000 198.240 346.100 200.240 ;
        RECT 4.000 196.840 345.700 198.240 ;
        RECT 4.000 188.040 346.100 196.840 ;
        RECT 4.400 186.640 346.100 188.040 ;
        RECT 4.000 184.640 346.100 186.640 ;
        RECT 4.000 183.240 345.700 184.640 ;
        RECT 4.000 174.440 346.100 183.240 ;
        RECT 4.400 173.040 346.100 174.440 ;
        RECT 4.000 171.040 346.100 173.040 ;
        RECT 4.000 169.640 345.700 171.040 ;
        RECT 4.000 160.840 346.100 169.640 ;
        RECT 4.400 159.440 346.100 160.840 ;
        RECT 4.000 157.440 346.100 159.440 ;
        RECT 4.000 156.040 345.700 157.440 ;
        RECT 4.000 147.240 346.100 156.040 ;
        RECT 4.400 145.840 346.100 147.240 ;
        RECT 4.000 143.840 346.100 145.840 ;
        RECT 4.000 142.440 345.700 143.840 ;
        RECT 4.000 133.640 346.100 142.440 ;
        RECT 4.400 132.240 346.100 133.640 ;
        RECT 4.000 130.240 346.100 132.240 ;
        RECT 4.000 128.840 345.700 130.240 ;
        RECT 4.000 120.040 346.100 128.840 ;
        RECT 4.400 118.640 346.100 120.040 ;
        RECT 4.000 116.640 346.100 118.640 ;
        RECT 4.000 115.240 345.700 116.640 ;
        RECT 4.000 106.440 346.100 115.240 ;
        RECT 4.400 105.040 346.100 106.440 ;
        RECT 4.000 103.040 346.100 105.040 ;
        RECT 4.000 101.640 345.700 103.040 ;
        RECT 4.000 92.840 346.100 101.640 ;
        RECT 4.400 91.440 346.100 92.840 ;
        RECT 4.000 89.440 346.100 91.440 ;
        RECT 4.000 88.040 345.700 89.440 ;
        RECT 4.000 79.240 346.100 88.040 ;
        RECT 4.400 77.840 346.100 79.240 ;
        RECT 4.000 75.840 346.100 77.840 ;
        RECT 4.000 74.440 345.700 75.840 ;
        RECT 4.000 65.640 346.100 74.440 ;
        RECT 4.400 64.240 346.100 65.640 ;
        RECT 4.000 62.240 346.100 64.240 ;
        RECT 4.000 60.840 345.700 62.240 ;
        RECT 4.000 52.040 346.100 60.840 ;
        RECT 4.400 50.640 346.100 52.040 ;
        RECT 4.000 48.640 346.100 50.640 ;
        RECT 4.000 47.240 345.700 48.640 ;
        RECT 4.000 38.440 346.100 47.240 ;
        RECT 4.400 37.040 346.100 38.440 ;
        RECT 4.000 35.040 346.100 37.040 ;
        RECT 4.000 33.640 345.700 35.040 ;
        RECT 4.000 24.840 346.100 33.640 ;
        RECT 4.400 23.440 346.100 24.840 ;
        RECT 4.000 21.440 346.100 23.440 ;
        RECT 4.000 20.040 345.700 21.440 ;
        RECT 4.000 11.240 346.100 20.040 ;
        RECT 4.400 9.840 346.100 11.240 ;
        RECT 4.000 7.840 346.100 9.840 ;
        RECT 4.000 6.975 345.700 7.840 ;
      LAYER met4 ;
        RECT 75.735 11.735 97.440 343.905 ;
        RECT 99.840 11.735 174.240 343.905 ;
        RECT 176.640 11.735 251.040 343.905 ;
        RECT 253.440 11.735 327.840 343.905 ;
        RECT 330.240 11.735 330.905 343.905 ;
  END
END wbuart_wrap
END LIBRARY

