magic
tech sky130A
magscale 1 2
timestamp 1654713014
<< obsli1 >>
rect 1104 2159 129720 130577
<< obsm1 >>
rect 290 144 130810 131232
<< metal2 >>
rect 386 132223 442 133023
rect 1122 132223 1178 133023
rect 1858 132223 1914 133023
rect 2686 132223 2742 133023
rect 3422 132223 3478 133023
rect 4250 132223 4306 133023
rect 4986 132223 5042 133023
rect 5722 132223 5778 133023
rect 6550 132223 6606 133023
rect 7286 132223 7342 133023
rect 8114 132223 8170 133023
rect 8850 132223 8906 133023
rect 9678 132223 9734 133023
rect 10414 132223 10470 133023
rect 11150 132223 11206 133023
rect 11978 132223 12034 133023
rect 12714 132223 12770 133023
rect 13542 132223 13598 133023
rect 14278 132223 14334 133023
rect 15014 132223 15070 133023
rect 15842 132223 15898 133023
rect 16578 132223 16634 133023
rect 17406 132223 17462 133023
rect 18142 132223 18198 133023
rect 18970 132223 19026 133023
rect 19706 132223 19762 133023
rect 20442 132223 20498 133023
rect 21270 132223 21326 133023
rect 22006 132223 22062 133023
rect 22834 132223 22890 133023
rect 23570 132223 23626 133023
rect 24398 132223 24454 133023
rect 25134 132223 25190 133023
rect 25870 132223 25926 133023
rect 26698 132223 26754 133023
rect 27434 132223 27490 133023
rect 28262 132223 28318 133023
rect 28998 132223 29054 133023
rect 29734 132223 29790 133023
rect 30562 132223 30618 133023
rect 31298 132223 31354 133023
rect 32126 132223 32182 133023
rect 32862 132223 32918 133023
rect 33690 132223 33746 133023
rect 34426 132223 34482 133023
rect 35162 132223 35218 133023
rect 35990 132223 36046 133023
rect 36726 132223 36782 133023
rect 37554 132223 37610 133023
rect 38290 132223 38346 133023
rect 39118 132223 39174 133023
rect 39854 132223 39910 133023
rect 40590 132223 40646 133023
rect 41418 132223 41474 133023
rect 42154 132223 42210 133023
rect 42982 132223 43038 133023
rect 43718 132223 43774 133023
rect 44454 132223 44510 133023
rect 45282 132223 45338 133023
rect 46018 132223 46074 133023
rect 46846 132223 46902 133023
rect 47582 132223 47638 133023
rect 48410 132223 48466 133023
rect 49146 132223 49202 133023
rect 49882 132223 49938 133023
rect 50710 132223 50766 133023
rect 51446 132223 51502 133023
rect 52274 132223 52330 133023
rect 53010 132223 53066 133023
rect 53746 132223 53802 133023
rect 54574 132223 54630 133023
rect 55310 132223 55366 133023
rect 56138 132223 56194 133023
rect 56874 132223 56930 133023
rect 57702 132223 57758 133023
rect 58438 132223 58494 133023
rect 59174 132223 59230 133023
rect 60002 132223 60058 133023
rect 60738 132223 60794 133023
rect 61566 132223 61622 133023
rect 62302 132223 62358 133023
rect 63130 132223 63186 133023
rect 63866 132223 63922 133023
rect 64602 132223 64658 133023
rect 65430 132223 65486 133023
rect 66166 132223 66222 133023
rect 66994 132223 67050 133023
rect 67730 132223 67786 133023
rect 68466 132223 68522 133023
rect 69294 132223 69350 133023
rect 70030 132223 70086 133023
rect 70858 132223 70914 133023
rect 71594 132223 71650 133023
rect 72422 132223 72478 133023
rect 73158 132223 73214 133023
rect 73894 132223 73950 133023
rect 74722 132223 74778 133023
rect 75458 132223 75514 133023
rect 76286 132223 76342 133023
rect 77022 132223 77078 133023
rect 77850 132223 77906 133023
rect 78586 132223 78642 133023
rect 79322 132223 79378 133023
rect 80150 132223 80206 133023
rect 80886 132223 80942 133023
rect 81714 132223 81770 133023
rect 82450 132223 82506 133023
rect 83186 132223 83242 133023
rect 84014 132223 84070 133023
rect 84750 132223 84806 133023
rect 85578 132223 85634 133023
rect 86314 132223 86370 133023
rect 87142 132223 87198 133023
rect 87878 132223 87934 133023
rect 88614 132223 88670 133023
rect 89442 132223 89498 133023
rect 90178 132223 90234 133023
rect 91006 132223 91062 133023
rect 91742 132223 91798 133023
rect 92478 132223 92534 133023
rect 93306 132223 93362 133023
rect 94042 132223 94098 133023
rect 94870 132223 94926 133023
rect 95606 132223 95662 133023
rect 96434 132223 96490 133023
rect 97170 132223 97226 133023
rect 97906 132223 97962 133023
rect 98734 132223 98790 133023
rect 99470 132223 99526 133023
rect 100298 132223 100354 133023
rect 101034 132223 101090 133023
rect 101862 132223 101918 133023
rect 102598 132223 102654 133023
rect 103334 132223 103390 133023
rect 104162 132223 104218 133023
rect 104898 132223 104954 133023
rect 105726 132223 105782 133023
rect 106462 132223 106518 133023
rect 107198 132223 107254 133023
rect 108026 132223 108082 133023
rect 108762 132223 108818 133023
rect 109590 132223 109646 133023
rect 110326 132223 110382 133023
rect 111154 132223 111210 133023
rect 111890 132223 111946 133023
rect 112626 132223 112682 133023
rect 113454 132223 113510 133023
rect 114190 132223 114246 133023
rect 115018 132223 115074 133023
rect 115754 132223 115810 133023
rect 116582 132223 116638 133023
rect 117318 132223 117374 133023
rect 118054 132223 118110 133023
rect 118882 132223 118938 133023
rect 119618 132223 119674 133023
rect 120446 132223 120502 133023
rect 121182 132223 121238 133023
rect 121918 132223 121974 133023
rect 122746 132223 122802 133023
rect 123482 132223 123538 133023
rect 124310 132223 124366 133023
rect 125046 132223 125102 133023
rect 125874 132223 125930 133023
rect 126610 132223 126666 133023
rect 127346 132223 127402 133023
rect 128174 132223 128230 133023
rect 128910 132223 128966 133023
rect 129738 132223 129794 133023
rect 130474 132223 130530 133023
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 754 0 810 800
rect 938 0 994 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5262 0 5318 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10690 0 10746 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16578 0 16634 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46754 0 46810 800
rect 46938 0 46994 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62578 0 62634 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63866 0 63922 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66074 0 66130 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67546 0 67602 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68650 0 68706 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 69938 0 69994 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70858 0 70914 800
rect 71042 0 71098 800
rect 71318 0 71374 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71962 0 72018 800
rect 72146 0 72202 800
rect 72330 0 72386 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73250 0 73306 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74538 0 74594 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75366 0 75422 800
rect 75642 0 75698 800
rect 75826 0 75882 800
rect 76010 0 76066 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80426 0 80482 800
rect 80610 0 80666 800
rect 80794 0 80850 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87602 0 87658 800
rect 87786 0 87842 800
rect 87970 0 88026 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90178 0 90234 800
rect 90362 0 90418 800
rect 90638 0 90694 800
rect 90822 0 90878 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91466 0 91522 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93674 0 93730 800
rect 93858 0 93914 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94502 0 94558 800
rect 94686 0 94742 800
rect 94962 0 95018 800
rect 95146 0 95202 800
rect 95330 0 95386 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97078 0 97134 800
rect 97354 0 97410 800
rect 97538 0 97594 800
rect 97722 0 97778 800
rect 97998 0 98054 800
rect 98182 0 98238 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99746 0 99802 800
rect 99930 0 99986 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100574 0 100630 800
rect 100758 0 100814 800
rect 101034 0 101090 800
rect 101218 0 101274 800
rect 101494 0 101550 800
rect 101678 0 101734 800
rect 101862 0 101918 800
rect 102138 0 102194 800
rect 102322 0 102378 800
rect 102506 0 102562 800
rect 102782 0 102838 800
rect 102966 0 103022 800
rect 103150 0 103206 800
rect 103426 0 103482 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104070 0 104126 800
rect 104254 0 104310 800
rect 104530 0 104586 800
rect 104714 0 104770 800
rect 104898 0 104954 800
rect 105174 0 105230 800
rect 105358 0 105414 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106002 0 106058 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106646 0 106702 800
rect 106922 0 106978 800
rect 107106 0 107162 800
rect 107290 0 107346 800
rect 107566 0 107622 800
rect 107750 0 107806 800
rect 107934 0 107990 800
rect 108210 0 108266 800
rect 108394 0 108450 800
rect 108578 0 108634 800
rect 108854 0 108910 800
rect 109038 0 109094 800
rect 109314 0 109370 800
rect 109498 0 109554 800
rect 109682 0 109738 800
rect 109958 0 110014 800
rect 110142 0 110198 800
rect 110326 0 110382 800
rect 110602 0 110658 800
rect 110786 0 110842 800
rect 110970 0 111026 800
rect 111246 0 111302 800
rect 111430 0 111486 800
rect 111614 0 111670 800
rect 111890 0 111946 800
rect 112074 0 112130 800
rect 112350 0 112406 800
rect 112534 0 112590 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113178 0 113234 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 113822 0 113878 800
rect 114006 0 114062 800
rect 114282 0 114338 800
rect 114466 0 114522 800
rect 114742 0 114798 800
rect 114926 0 114982 800
rect 115110 0 115166 800
rect 115386 0 115442 800
rect 115570 0 115626 800
rect 115754 0 115810 800
rect 116030 0 116086 800
rect 116214 0 116270 800
rect 116398 0 116454 800
rect 116674 0 116730 800
rect 116858 0 116914 800
rect 117042 0 117098 800
rect 117318 0 117374 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 117962 0 118018 800
rect 118146 0 118202 800
rect 118422 0 118478 800
rect 118606 0 118662 800
rect 118790 0 118846 800
rect 119066 0 119122 800
rect 119250 0 119306 800
rect 119434 0 119490 800
rect 119710 0 119766 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120354 0 120410 800
rect 120538 0 120594 800
rect 120814 0 120870 800
rect 120998 0 121054 800
rect 121182 0 121238 800
rect 121458 0 121514 800
rect 121642 0 121698 800
rect 121826 0 121882 800
rect 122102 0 122158 800
rect 122286 0 122342 800
rect 122470 0 122526 800
rect 122746 0 122802 800
rect 122930 0 122986 800
rect 123206 0 123262 800
rect 123390 0 123446 800
rect 123574 0 123630 800
rect 123850 0 123906 800
rect 124034 0 124090 800
rect 124218 0 124274 800
rect 124494 0 124550 800
rect 124678 0 124734 800
rect 124862 0 124918 800
rect 125138 0 125194 800
rect 125322 0 125378 800
rect 125598 0 125654 800
rect 125782 0 125838 800
rect 125966 0 126022 800
rect 126242 0 126298 800
rect 126426 0 126482 800
rect 126610 0 126666 800
rect 126886 0 126942 800
rect 127070 0 127126 800
rect 127254 0 127310 800
rect 127530 0 127586 800
rect 127714 0 127770 800
rect 127898 0 127954 800
rect 128174 0 128230 800
rect 128358 0 128414 800
rect 128634 0 128690 800
rect 128818 0 128874 800
rect 129002 0 129058 800
rect 129278 0 129334 800
rect 129462 0 129518 800
rect 129646 0 129702 800
rect 129922 0 129978 800
rect 130106 0 130162 800
rect 130290 0 130346 800
rect 130566 0 130622 800
rect 130750 0 130806 800
<< obsm2 >>
rect 18 132167 330 132274
rect 498 132167 1066 132274
rect 1234 132167 1802 132274
rect 1970 132167 2630 132274
rect 2798 132167 3366 132274
rect 3534 132167 4194 132274
rect 4362 132167 4930 132274
rect 5098 132167 5666 132274
rect 5834 132167 6494 132274
rect 6662 132167 7230 132274
rect 7398 132167 8058 132274
rect 8226 132167 8794 132274
rect 8962 132167 9622 132274
rect 9790 132167 10358 132274
rect 10526 132167 11094 132274
rect 11262 132167 11922 132274
rect 12090 132167 12658 132274
rect 12826 132167 13486 132274
rect 13654 132167 14222 132274
rect 14390 132167 14958 132274
rect 15126 132167 15786 132274
rect 15954 132167 16522 132274
rect 16690 132167 17350 132274
rect 17518 132167 18086 132274
rect 18254 132167 18914 132274
rect 19082 132167 19650 132274
rect 19818 132167 20386 132274
rect 20554 132167 21214 132274
rect 21382 132167 21950 132274
rect 22118 132167 22778 132274
rect 22946 132167 23514 132274
rect 23682 132167 24342 132274
rect 24510 132167 25078 132274
rect 25246 132167 25814 132274
rect 25982 132167 26642 132274
rect 26810 132167 27378 132274
rect 27546 132167 28206 132274
rect 28374 132167 28942 132274
rect 29110 132167 29678 132274
rect 29846 132167 30506 132274
rect 30674 132167 31242 132274
rect 31410 132167 32070 132274
rect 32238 132167 32806 132274
rect 32974 132167 33634 132274
rect 33802 132167 34370 132274
rect 34538 132167 35106 132274
rect 35274 132167 35934 132274
rect 36102 132167 36670 132274
rect 36838 132167 37498 132274
rect 37666 132167 38234 132274
rect 38402 132167 39062 132274
rect 39230 132167 39798 132274
rect 39966 132167 40534 132274
rect 40702 132167 41362 132274
rect 41530 132167 42098 132274
rect 42266 132167 42926 132274
rect 43094 132167 43662 132274
rect 43830 132167 44398 132274
rect 44566 132167 45226 132274
rect 45394 132167 45962 132274
rect 46130 132167 46790 132274
rect 46958 132167 47526 132274
rect 47694 132167 48354 132274
rect 48522 132167 49090 132274
rect 49258 132167 49826 132274
rect 49994 132167 50654 132274
rect 50822 132167 51390 132274
rect 51558 132167 52218 132274
rect 52386 132167 52954 132274
rect 53122 132167 53690 132274
rect 53858 132167 54518 132274
rect 54686 132167 55254 132274
rect 55422 132167 56082 132274
rect 56250 132167 56818 132274
rect 56986 132167 57646 132274
rect 57814 132167 58382 132274
rect 58550 132167 59118 132274
rect 59286 132167 59946 132274
rect 60114 132167 60682 132274
rect 60850 132167 61510 132274
rect 61678 132167 62246 132274
rect 62414 132167 63074 132274
rect 63242 132167 63810 132274
rect 63978 132167 64546 132274
rect 64714 132167 65374 132274
rect 65542 132167 66110 132274
rect 66278 132167 66938 132274
rect 67106 132167 67674 132274
rect 67842 132167 68410 132274
rect 68578 132167 69238 132274
rect 69406 132167 69974 132274
rect 70142 132167 70802 132274
rect 70970 132167 71538 132274
rect 71706 132167 72366 132274
rect 72534 132167 73102 132274
rect 73270 132167 73838 132274
rect 74006 132167 74666 132274
rect 74834 132167 75402 132274
rect 75570 132167 76230 132274
rect 76398 132167 76966 132274
rect 77134 132167 77794 132274
rect 77962 132167 78530 132274
rect 78698 132167 79266 132274
rect 79434 132167 80094 132274
rect 80262 132167 80830 132274
rect 80998 132167 81658 132274
rect 81826 132167 82394 132274
rect 82562 132167 83130 132274
rect 83298 132167 83958 132274
rect 84126 132167 84694 132274
rect 84862 132167 85522 132274
rect 85690 132167 86258 132274
rect 86426 132167 87086 132274
rect 87254 132167 87822 132274
rect 87990 132167 88558 132274
rect 88726 132167 89386 132274
rect 89554 132167 90122 132274
rect 90290 132167 90950 132274
rect 91118 132167 91686 132274
rect 91854 132167 92422 132274
rect 92590 132167 93250 132274
rect 93418 132167 93986 132274
rect 94154 132167 94814 132274
rect 94982 132167 95550 132274
rect 95718 132167 96378 132274
rect 96546 132167 97114 132274
rect 97282 132167 97850 132274
rect 98018 132167 98678 132274
rect 98846 132167 99414 132274
rect 99582 132167 100242 132274
rect 100410 132167 100978 132274
rect 101146 132167 101806 132274
rect 101974 132167 102542 132274
rect 102710 132167 103278 132274
rect 103446 132167 104106 132274
rect 104274 132167 104842 132274
rect 105010 132167 105670 132274
rect 105838 132167 106406 132274
rect 106574 132167 107142 132274
rect 107310 132167 107970 132274
rect 108138 132167 108706 132274
rect 108874 132167 109534 132274
rect 109702 132167 110270 132274
rect 110438 132167 111098 132274
rect 111266 132167 111834 132274
rect 112002 132167 112570 132274
rect 112738 132167 113398 132274
rect 113566 132167 114134 132274
rect 114302 132167 114962 132274
rect 115130 132167 115698 132274
rect 115866 132167 116526 132274
rect 116694 132167 117262 132274
rect 117430 132167 117998 132274
rect 118166 132167 118826 132274
rect 118994 132167 119562 132274
rect 119730 132167 120390 132274
rect 120558 132167 121126 132274
rect 121294 132167 121862 132274
rect 122030 132167 122690 132274
rect 122858 132167 123426 132274
rect 123594 132167 124254 132274
rect 124422 132167 124990 132274
rect 125158 132167 125818 132274
rect 125986 132167 126554 132274
rect 126722 132167 127290 132274
rect 127458 132167 128118 132274
rect 128286 132167 128854 132274
rect 129022 132167 129682 132274
rect 129850 132167 130418 132274
rect 130586 132167 130804 132274
rect 18 856 130804 132167
rect 18 138 54 856
rect 222 138 238 856
rect 406 138 422 856
rect 590 138 698 856
rect 866 138 882 856
rect 1050 138 1066 856
rect 1234 138 1342 856
rect 1510 138 1526 856
rect 1694 138 1710 856
rect 1878 138 1986 856
rect 2154 138 2170 856
rect 2338 138 2354 856
rect 2522 138 2630 856
rect 2798 138 2814 856
rect 2982 138 3090 856
rect 3258 138 3274 856
rect 3442 138 3458 856
rect 3626 138 3734 856
rect 3902 138 3918 856
rect 4086 138 4102 856
rect 4270 138 4378 856
rect 4546 138 4562 856
rect 4730 138 4746 856
rect 4914 138 5022 856
rect 5190 138 5206 856
rect 5374 138 5390 856
rect 5558 138 5666 856
rect 5834 138 5850 856
rect 6018 138 6126 856
rect 6294 138 6310 856
rect 6478 138 6494 856
rect 6662 138 6770 856
rect 6938 138 6954 856
rect 7122 138 7138 856
rect 7306 138 7414 856
rect 7582 138 7598 856
rect 7766 138 7782 856
rect 7950 138 8058 856
rect 8226 138 8242 856
rect 8410 138 8518 856
rect 8686 138 8702 856
rect 8870 138 8886 856
rect 9054 138 9162 856
rect 9330 138 9346 856
rect 9514 138 9530 856
rect 9698 138 9806 856
rect 9974 138 9990 856
rect 10158 138 10174 856
rect 10342 138 10450 856
rect 10618 138 10634 856
rect 10802 138 10818 856
rect 10986 138 11094 856
rect 11262 138 11278 856
rect 11446 138 11554 856
rect 11722 138 11738 856
rect 11906 138 11922 856
rect 12090 138 12198 856
rect 12366 138 12382 856
rect 12550 138 12566 856
rect 12734 138 12842 856
rect 13010 138 13026 856
rect 13194 138 13210 856
rect 13378 138 13486 856
rect 13654 138 13670 856
rect 13838 138 13946 856
rect 14114 138 14130 856
rect 14298 138 14314 856
rect 14482 138 14590 856
rect 14758 138 14774 856
rect 14942 138 14958 856
rect 15126 138 15234 856
rect 15402 138 15418 856
rect 15586 138 15602 856
rect 15770 138 15878 856
rect 16046 138 16062 856
rect 16230 138 16246 856
rect 16414 138 16522 856
rect 16690 138 16706 856
rect 16874 138 16982 856
rect 17150 138 17166 856
rect 17334 138 17350 856
rect 17518 138 17626 856
rect 17794 138 17810 856
rect 17978 138 17994 856
rect 18162 138 18270 856
rect 18438 138 18454 856
rect 18622 138 18638 856
rect 18806 138 18914 856
rect 19082 138 19098 856
rect 19266 138 19374 856
rect 19542 138 19558 856
rect 19726 138 19742 856
rect 19910 138 20018 856
rect 20186 138 20202 856
rect 20370 138 20386 856
rect 20554 138 20662 856
rect 20830 138 20846 856
rect 21014 138 21030 856
rect 21198 138 21306 856
rect 21474 138 21490 856
rect 21658 138 21674 856
rect 21842 138 21950 856
rect 22118 138 22134 856
rect 22302 138 22410 856
rect 22578 138 22594 856
rect 22762 138 22778 856
rect 22946 138 23054 856
rect 23222 138 23238 856
rect 23406 138 23422 856
rect 23590 138 23698 856
rect 23866 138 23882 856
rect 24050 138 24066 856
rect 24234 138 24342 856
rect 24510 138 24526 856
rect 24694 138 24802 856
rect 24970 138 24986 856
rect 25154 138 25170 856
rect 25338 138 25446 856
rect 25614 138 25630 856
rect 25798 138 25814 856
rect 25982 138 26090 856
rect 26258 138 26274 856
rect 26442 138 26458 856
rect 26626 138 26734 856
rect 26902 138 26918 856
rect 27086 138 27102 856
rect 27270 138 27378 856
rect 27546 138 27562 856
rect 27730 138 27838 856
rect 28006 138 28022 856
rect 28190 138 28206 856
rect 28374 138 28482 856
rect 28650 138 28666 856
rect 28834 138 28850 856
rect 29018 138 29126 856
rect 29294 138 29310 856
rect 29478 138 29494 856
rect 29662 138 29770 856
rect 29938 138 29954 856
rect 30122 138 30230 856
rect 30398 138 30414 856
rect 30582 138 30598 856
rect 30766 138 30874 856
rect 31042 138 31058 856
rect 31226 138 31242 856
rect 31410 138 31518 856
rect 31686 138 31702 856
rect 31870 138 31886 856
rect 32054 138 32162 856
rect 32330 138 32346 856
rect 32514 138 32530 856
rect 32698 138 32806 856
rect 32974 138 32990 856
rect 33158 138 33266 856
rect 33434 138 33450 856
rect 33618 138 33634 856
rect 33802 138 33910 856
rect 34078 138 34094 856
rect 34262 138 34278 856
rect 34446 138 34554 856
rect 34722 138 34738 856
rect 34906 138 34922 856
rect 35090 138 35198 856
rect 35366 138 35382 856
rect 35550 138 35658 856
rect 35826 138 35842 856
rect 36010 138 36026 856
rect 36194 138 36302 856
rect 36470 138 36486 856
rect 36654 138 36670 856
rect 36838 138 36946 856
rect 37114 138 37130 856
rect 37298 138 37314 856
rect 37482 138 37590 856
rect 37758 138 37774 856
rect 37942 138 37958 856
rect 38126 138 38234 856
rect 38402 138 38418 856
rect 38586 138 38694 856
rect 38862 138 38878 856
rect 39046 138 39062 856
rect 39230 138 39338 856
rect 39506 138 39522 856
rect 39690 138 39706 856
rect 39874 138 39982 856
rect 40150 138 40166 856
rect 40334 138 40350 856
rect 40518 138 40626 856
rect 40794 138 40810 856
rect 40978 138 41086 856
rect 41254 138 41270 856
rect 41438 138 41454 856
rect 41622 138 41730 856
rect 41898 138 41914 856
rect 42082 138 42098 856
rect 42266 138 42374 856
rect 42542 138 42558 856
rect 42726 138 42742 856
rect 42910 138 43018 856
rect 43186 138 43202 856
rect 43370 138 43386 856
rect 43554 138 43662 856
rect 43830 138 43846 856
rect 44014 138 44122 856
rect 44290 138 44306 856
rect 44474 138 44490 856
rect 44658 138 44766 856
rect 44934 138 44950 856
rect 45118 138 45134 856
rect 45302 138 45410 856
rect 45578 138 45594 856
rect 45762 138 45778 856
rect 45946 138 46054 856
rect 46222 138 46238 856
rect 46406 138 46514 856
rect 46682 138 46698 856
rect 46866 138 46882 856
rect 47050 138 47158 856
rect 47326 138 47342 856
rect 47510 138 47526 856
rect 47694 138 47802 856
rect 47970 138 47986 856
rect 48154 138 48170 856
rect 48338 138 48446 856
rect 48614 138 48630 856
rect 48798 138 48814 856
rect 48982 138 49090 856
rect 49258 138 49274 856
rect 49442 138 49550 856
rect 49718 138 49734 856
rect 49902 138 49918 856
rect 50086 138 50194 856
rect 50362 138 50378 856
rect 50546 138 50562 856
rect 50730 138 50838 856
rect 51006 138 51022 856
rect 51190 138 51206 856
rect 51374 138 51482 856
rect 51650 138 51666 856
rect 51834 138 51942 856
rect 52110 138 52126 856
rect 52294 138 52310 856
rect 52478 138 52586 856
rect 52754 138 52770 856
rect 52938 138 52954 856
rect 53122 138 53230 856
rect 53398 138 53414 856
rect 53582 138 53598 856
rect 53766 138 53874 856
rect 54042 138 54058 856
rect 54226 138 54242 856
rect 54410 138 54518 856
rect 54686 138 54702 856
rect 54870 138 54978 856
rect 55146 138 55162 856
rect 55330 138 55346 856
rect 55514 138 55622 856
rect 55790 138 55806 856
rect 55974 138 55990 856
rect 56158 138 56266 856
rect 56434 138 56450 856
rect 56618 138 56634 856
rect 56802 138 56910 856
rect 57078 138 57094 856
rect 57262 138 57370 856
rect 57538 138 57554 856
rect 57722 138 57738 856
rect 57906 138 58014 856
rect 58182 138 58198 856
rect 58366 138 58382 856
rect 58550 138 58658 856
rect 58826 138 58842 856
rect 59010 138 59026 856
rect 59194 138 59302 856
rect 59470 138 59486 856
rect 59654 138 59670 856
rect 59838 138 59946 856
rect 60114 138 60130 856
rect 60298 138 60406 856
rect 60574 138 60590 856
rect 60758 138 60774 856
rect 60942 138 61050 856
rect 61218 138 61234 856
rect 61402 138 61418 856
rect 61586 138 61694 856
rect 61862 138 61878 856
rect 62046 138 62062 856
rect 62230 138 62338 856
rect 62506 138 62522 856
rect 62690 138 62798 856
rect 62966 138 62982 856
rect 63150 138 63166 856
rect 63334 138 63442 856
rect 63610 138 63626 856
rect 63794 138 63810 856
rect 63978 138 64086 856
rect 64254 138 64270 856
rect 64438 138 64454 856
rect 64622 138 64730 856
rect 64898 138 64914 856
rect 65082 138 65098 856
rect 65266 138 65374 856
rect 65542 138 65558 856
rect 65726 138 65834 856
rect 66002 138 66018 856
rect 66186 138 66202 856
rect 66370 138 66478 856
rect 66646 138 66662 856
rect 66830 138 66846 856
rect 67014 138 67122 856
rect 67290 138 67306 856
rect 67474 138 67490 856
rect 67658 138 67766 856
rect 67934 138 67950 856
rect 68118 138 68134 856
rect 68302 138 68410 856
rect 68578 138 68594 856
rect 68762 138 68870 856
rect 69038 138 69054 856
rect 69222 138 69238 856
rect 69406 138 69514 856
rect 69682 138 69698 856
rect 69866 138 69882 856
rect 70050 138 70158 856
rect 70326 138 70342 856
rect 70510 138 70526 856
rect 70694 138 70802 856
rect 70970 138 70986 856
rect 71154 138 71262 856
rect 71430 138 71446 856
rect 71614 138 71630 856
rect 71798 138 71906 856
rect 72074 138 72090 856
rect 72258 138 72274 856
rect 72442 138 72550 856
rect 72718 138 72734 856
rect 72902 138 72918 856
rect 73086 138 73194 856
rect 73362 138 73378 856
rect 73546 138 73562 856
rect 73730 138 73838 856
rect 74006 138 74022 856
rect 74190 138 74298 856
rect 74466 138 74482 856
rect 74650 138 74666 856
rect 74834 138 74942 856
rect 75110 138 75126 856
rect 75294 138 75310 856
rect 75478 138 75586 856
rect 75754 138 75770 856
rect 75938 138 75954 856
rect 76122 138 76230 856
rect 76398 138 76414 856
rect 76582 138 76690 856
rect 76858 138 76874 856
rect 77042 138 77058 856
rect 77226 138 77334 856
rect 77502 138 77518 856
rect 77686 138 77702 856
rect 77870 138 77978 856
rect 78146 138 78162 856
rect 78330 138 78346 856
rect 78514 138 78622 856
rect 78790 138 78806 856
rect 78974 138 78990 856
rect 79158 138 79266 856
rect 79434 138 79450 856
rect 79618 138 79726 856
rect 79894 138 79910 856
rect 80078 138 80094 856
rect 80262 138 80370 856
rect 80538 138 80554 856
rect 80722 138 80738 856
rect 80906 138 81014 856
rect 81182 138 81198 856
rect 81366 138 81382 856
rect 81550 138 81658 856
rect 81826 138 81842 856
rect 82010 138 82118 856
rect 82286 138 82302 856
rect 82470 138 82486 856
rect 82654 138 82762 856
rect 82930 138 82946 856
rect 83114 138 83130 856
rect 83298 138 83406 856
rect 83574 138 83590 856
rect 83758 138 83774 856
rect 83942 138 84050 856
rect 84218 138 84234 856
rect 84402 138 84418 856
rect 84586 138 84694 856
rect 84862 138 84878 856
rect 85046 138 85154 856
rect 85322 138 85338 856
rect 85506 138 85522 856
rect 85690 138 85798 856
rect 85966 138 85982 856
rect 86150 138 86166 856
rect 86334 138 86442 856
rect 86610 138 86626 856
rect 86794 138 86810 856
rect 86978 138 87086 856
rect 87254 138 87270 856
rect 87438 138 87546 856
rect 87714 138 87730 856
rect 87898 138 87914 856
rect 88082 138 88190 856
rect 88358 138 88374 856
rect 88542 138 88558 856
rect 88726 138 88834 856
rect 89002 138 89018 856
rect 89186 138 89202 856
rect 89370 138 89478 856
rect 89646 138 89662 856
rect 89830 138 89846 856
rect 90014 138 90122 856
rect 90290 138 90306 856
rect 90474 138 90582 856
rect 90750 138 90766 856
rect 90934 138 90950 856
rect 91118 138 91226 856
rect 91394 138 91410 856
rect 91578 138 91594 856
rect 91762 138 91870 856
rect 92038 138 92054 856
rect 92222 138 92238 856
rect 92406 138 92514 856
rect 92682 138 92698 856
rect 92866 138 92974 856
rect 93142 138 93158 856
rect 93326 138 93342 856
rect 93510 138 93618 856
rect 93786 138 93802 856
rect 93970 138 93986 856
rect 94154 138 94262 856
rect 94430 138 94446 856
rect 94614 138 94630 856
rect 94798 138 94906 856
rect 95074 138 95090 856
rect 95258 138 95274 856
rect 95442 138 95550 856
rect 95718 138 95734 856
rect 95902 138 96010 856
rect 96178 138 96194 856
rect 96362 138 96378 856
rect 96546 138 96654 856
rect 96822 138 96838 856
rect 97006 138 97022 856
rect 97190 138 97298 856
rect 97466 138 97482 856
rect 97650 138 97666 856
rect 97834 138 97942 856
rect 98110 138 98126 856
rect 98294 138 98402 856
rect 98570 138 98586 856
rect 98754 138 98770 856
rect 98938 138 99046 856
rect 99214 138 99230 856
rect 99398 138 99414 856
rect 99582 138 99690 856
rect 99858 138 99874 856
rect 100042 138 100058 856
rect 100226 138 100334 856
rect 100502 138 100518 856
rect 100686 138 100702 856
rect 100870 138 100978 856
rect 101146 138 101162 856
rect 101330 138 101438 856
rect 101606 138 101622 856
rect 101790 138 101806 856
rect 101974 138 102082 856
rect 102250 138 102266 856
rect 102434 138 102450 856
rect 102618 138 102726 856
rect 102894 138 102910 856
rect 103078 138 103094 856
rect 103262 138 103370 856
rect 103538 138 103554 856
rect 103722 138 103830 856
rect 103998 138 104014 856
rect 104182 138 104198 856
rect 104366 138 104474 856
rect 104642 138 104658 856
rect 104826 138 104842 856
rect 105010 138 105118 856
rect 105286 138 105302 856
rect 105470 138 105486 856
rect 105654 138 105762 856
rect 105930 138 105946 856
rect 106114 138 106130 856
rect 106298 138 106406 856
rect 106574 138 106590 856
rect 106758 138 106866 856
rect 107034 138 107050 856
rect 107218 138 107234 856
rect 107402 138 107510 856
rect 107678 138 107694 856
rect 107862 138 107878 856
rect 108046 138 108154 856
rect 108322 138 108338 856
rect 108506 138 108522 856
rect 108690 138 108798 856
rect 108966 138 108982 856
rect 109150 138 109258 856
rect 109426 138 109442 856
rect 109610 138 109626 856
rect 109794 138 109902 856
rect 110070 138 110086 856
rect 110254 138 110270 856
rect 110438 138 110546 856
rect 110714 138 110730 856
rect 110898 138 110914 856
rect 111082 138 111190 856
rect 111358 138 111374 856
rect 111542 138 111558 856
rect 111726 138 111834 856
rect 112002 138 112018 856
rect 112186 138 112294 856
rect 112462 138 112478 856
rect 112646 138 112662 856
rect 112830 138 112938 856
rect 113106 138 113122 856
rect 113290 138 113306 856
rect 113474 138 113582 856
rect 113750 138 113766 856
rect 113934 138 113950 856
rect 114118 138 114226 856
rect 114394 138 114410 856
rect 114578 138 114686 856
rect 114854 138 114870 856
rect 115038 138 115054 856
rect 115222 138 115330 856
rect 115498 138 115514 856
rect 115682 138 115698 856
rect 115866 138 115974 856
rect 116142 138 116158 856
rect 116326 138 116342 856
rect 116510 138 116618 856
rect 116786 138 116802 856
rect 116970 138 116986 856
rect 117154 138 117262 856
rect 117430 138 117446 856
rect 117614 138 117722 856
rect 117890 138 117906 856
rect 118074 138 118090 856
rect 118258 138 118366 856
rect 118534 138 118550 856
rect 118718 138 118734 856
rect 118902 138 119010 856
rect 119178 138 119194 856
rect 119362 138 119378 856
rect 119546 138 119654 856
rect 119822 138 119838 856
rect 120006 138 120114 856
rect 120282 138 120298 856
rect 120466 138 120482 856
rect 120650 138 120758 856
rect 120926 138 120942 856
rect 121110 138 121126 856
rect 121294 138 121402 856
rect 121570 138 121586 856
rect 121754 138 121770 856
rect 121938 138 122046 856
rect 122214 138 122230 856
rect 122398 138 122414 856
rect 122582 138 122690 856
rect 122858 138 122874 856
rect 123042 138 123150 856
rect 123318 138 123334 856
rect 123502 138 123518 856
rect 123686 138 123794 856
rect 123962 138 123978 856
rect 124146 138 124162 856
rect 124330 138 124438 856
rect 124606 138 124622 856
rect 124790 138 124806 856
rect 124974 138 125082 856
rect 125250 138 125266 856
rect 125434 138 125542 856
rect 125710 138 125726 856
rect 125894 138 125910 856
rect 126078 138 126186 856
rect 126354 138 126370 856
rect 126538 138 126554 856
rect 126722 138 126830 856
rect 126998 138 127014 856
rect 127182 138 127198 856
rect 127366 138 127474 856
rect 127642 138 127658 856
rect 127826 138 127842 856
rect 128010 138 128118 856
rect 128286 138 128302 856
rect 128470 138 128578 856
rect 128746 138 128762 856
rect 128930 138 128946 856
rect 129114 138 129222 856
rect 129390 138 129406 856
rect 129574 138 129590 856
rect 129758 138 129866 856
rect 130034 138 130050 856
rect 130218 138 130234 856
rect 130402 138 130510 856
rect 130678 138 130694 856
<< obsm3 >>
rect 13 307 128787 131069
<< metal4 >>
rect 4208 2128 4528 130608
rect 19568 2128 19888 130608
rect 34928 2128 35248 130608
rect 50288 2128 50608 130608
rect 65648 2128 65968 130608
rect 81008 2128 81328 130608
rect 96368 2128 96688 130608
rect 111728 2128 112048 130608
rect 127088 2128 127408 130608
<< obsm4 >>
rect 2083 130688 128189 131069
rect 2083 2048 4128 130688
rect 4608 2048 19488 130688
rect 19968 2048 34848 130688
rect 35328 2048 50208 130688
rect 50688 2048 65568 130688
rect 66048 2048 80928 130688
rect 81408 2048 96288 130688
rect 96768 2048 111648 130688
rect 112128 2048 127008 130688
rect 127488 2048 128189 130688
rect 2083 307 128189 2048
<< labels >>
rlabel metal2 s 2686 132223 2742 133023 6 dram_addr0[0]
port 1 nsew signal output
rlabel metal2 s 5722 132223 5778 133023 6 dram_addr0[1]
port 2 nsew signal output
rlabel metal2 s 8850 132223 8906 133023 6 dram_addr0[2]
port 3 nsew signal output
rlabel metal2 s 11978 132223 12034 133023 6 dram_addr0[3]
port 4 nsew signal output
rlabel metal2 s 15014 132223 15070 133023 6 dram_addr0[4]
port 5 nsew signal output
rlabel metal2 s 17406 132223 17462 133023 6 dram_addr0[5]
port 6 nsew signal output
rlabel metal2 s 19706 132223 19762 133023 6 dram_addr0[6]
port 7 nsew signal output
rlabel metal2 s 22006 132223 22062 133023 6 dram_addr0[7]
port 8 nsew signal output
rlabel metal2 s 24398 132223 24454 133023 6 dram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 386 132223 442 133023 6 dram_clk0
port 10 nsew signal output
rlabel metal2 s 1122 132223 1178 133023 6 dram_csb0
port 11 nsew signal output
rlabel metal2 s 3422 132223 3478 133023 6 dram_din0[0]
port 12 nsew signal output
rlabel metal2 s 28262 132223 28318 133023 6 dram_din0[10]
port 13 nsew signal output
rlabel metal2 s 29734 132223 29790 133023 6 dram_din0[11]
port 14 nsew signal output
rlabel metal2 s 31298 132223 31354 133023 6 dram_din0[12]
port 15 nsew signal output
rlabel metal2 s 32862 132223 32918 133023 6 dram_din0[13]
port 16 nsew signal output
rlabel metal2 s 34426 132223 34482 133023 6 dram_din0[14]
port 17 nsew signal output
rlabel metal2 s 35990 132223 36046 133023 6 dram_din0[15]
port 18 nsew signal output
rlabel metal2 s 37554 132223 37610 133023 6 dram_din0[16]
port 19 nsew signal output
rlabel metal2 s 39118 132223 39174 133023 6 dram_din0[17]
port 20 nsew signal output
rlabel metal2 s 40590 132223 40646 133023 6 dram_din0[18]
port 21 nsew signal output
rlabel metal2 s 42154 132223 42210 133023 6 dram_din0[19]
port 22 nsew signal output
rlabel metal2 s 6550 132223 6606 133023 6 dram_din0[1]
port 23 nsew signal output
rlabel metal2 s 43718 132223 43774 133023 6 dram_din0[20]
port 24 nsew signal output
rlabel metal2 s 45282 132223 45338 133023 6 dram_din0[21]
port 25 nsew signal output
rlabel metal2 s 46846 132223 46902 133023 6 dram_din0[22]
port 26 nsew signal output
rlabel metal2 s 48410 132223 48466 133023 6 dram_din0[23]
port 27 nsew signal output
rlabel metal2 s 49882 132223 49938 133023 6 dram_din0[24]
port 28 nsew signal output
rlabel metal2 s 51446 132223 51502 133023 6 dram_din0[25]
port 29 nsew signal output
rlabel metal2 s 53010 132223 53066 133023 6 dram_din0[26]
port 30 nsew signal output
rlabel metal2 s 54574 132223 54630 133023 6 dram_din0[27]
port 31 nsew signal output
rlabel metal2 s 56138 132223 56194 133023 6 dram_din0[28]
port 32 nsew signal output
rlabel metal2 s 57702 132223 57758 133023 6 dram_din0[29]
port 33 nsew signal output
rlabel metal2 s 9678 132223 9734 133023 6 dram_din0[2]
port 34 nsew signal output
rlabel metal2 s 59174 132223 59230 133023 6 dram_din0[30]
port 35 nsew signal output
rlabel metal2 s 60738 132223 60794 133023 6 dram_din0[31]
port 36 nsew signal output
rlabel metal2 s 12714 132223 12770 133023 6 dram_din0[3]
port 37 nsew signal output
rlabel metal2 s 15842 132223 15898 133023 6 dram_din0[4]
port 38 nsew signal output
rlabel metal2 s 18142 132223 18198 133023 6 dram_din0[5]
port 39 nsew signal output
rlabel metal2 s 20442 132223 20498 133023 6 dram_din0[6]
port 40 nsew signal output
rlabel metal2 s 22834 132223 22890 133023 6 dram_din0[7]
port 41 nsew signal output
rlabel metal2 s 25134 132223 25190 133023 6 dram_din0[8]
port 42 nsew signal output
rlabel metal2 s 26698 132223 26754 133023 6 dram_din0[9]
port 43 nsew signal output
rlabel metal2 s 4250 132223 4306 133023 6 dram_dout0[0]
port 44 nsew signal input
rlabel metal2 s 28998 132223 29054 133023 6 dram_dout0[10]
port 45 nsew signal input
rlabel metal2 s 30562 132223 30618 133023 6 dram_dout0[11]
port 46 nsew signal input
rlabel metal2 s 32126 132223 32182 133023 6 dram_dout0[12]
port 47 nsew signal input
rlabel metal2 s 33690 132223 33746 133023 6 dram_dout0[13]
port 48 nsew signal input
rlabel metal2 s 35162 132223 35218 133023 6 dram_dout0[14]
port 49 nsew signal input
rlabel metal2 s 36726 132223 36782 133023 6 dram_dout0[15]
port 50 nsew signal input
rlabel metal2 s 38290 132223 38346 133023 6 dram_dout0[16]
port 51 nsew signal input
rlabel metal2 s 39854 132223 39910 133023 6 dram_dout0[17]
port 52 nsew signal input
rlabel metal2 s 41418 132223 41474 133023 6 dram_dout0[18]
port 53 nsew signal input
rlabel metal2 s 42982 132223 43038 133023 6 dram_dout0[19]
port 54 nsew signal input
rlabel metal2 s 7286 132223 7342 133023 6 dram_dout0[1]
port 55 nsew signal input
rlabel metal2 s 44454 132223 44510 133023 6 dram_dout0[20]
port 56 nsew signal input
rlabel metal2 s 46018 132223 46074 133023 6 dram_dout0[21]
port 57 nsew signal input
rlabel metal2 s 47582 132223 47638 133023 6 dram_dout0[22]
port 58 nsew signal input
rlabel metal2 s 49146 132223 49202 133023 6 dram_dout0[23]
port 59 nsew signal input
rlabel metal2 s 50710 132223 50766 133023 6 dram_dout0[24]
port 60 nsew signal input
rlabel metal2 s 52274 132223 52330 133023 6 dram_dout0[25]
port 61 nsew signal input
rlabel metal2 s 53746 132223 53802 133023 6 dram_dout0[26]
port 62 nsew signal input
rlabel metal2 s 55310 132223 55366 133023 6 dram_dout0[27]
port 63 nsew signal input
rlabel metal2 s 56874 132223 56930 133023 6 dram_dout0[28]
port 64 nsew signal input
rlabel metal2 s 58438 132223 58494 133023 6 dram_dout0[29]
port 65 nsew signal input
rlabel metal2 s 10414 132223 10470 133023 6 dram_dout0[2]
port 66 nsew signal input
rlabel metal2 s 60002 132223 60058 133023 6 dram_dout0[30]
port 67 nsew signal input
rlabel metal2 s 61566 132223 61622 133023 6 dram_dout0[31]
port 68 nsew signal input
rlabel metal2 s 13542 132223 13598 133023 6 dram_dout0[3]
port 69 nsew signal input
rlabel metal2 s 16578 132223 16634 133023 6 dram_dout0[4]
port 70 nsew signal input
rlabel metal2 s 18970 132223 19026 133023 6 dram_dout0[5]
port 71 nsew signal input
rlabel metal2 s 21270 132223 21326 133023 6 dram_dout0[6]
port 72 nsew signal input
rlabel metal2 s 23570 132223 23626 133023 6 dram_dout0[7]
port 73 nsew signal input
rlabel metal2 s 25870 132223 25926 133023 6 dram_dout0[8]
port 74 nsew signal input
rlabel metal2 s 27434 132223 27490 133023 6 dram_dout0[9]
port 75 nsew signal input
rlabel metal2 s 1858 132223 1914 133023 6 dram_web0
port 76 nsew signal output
rlabel metal2 s 4986 132223 5042 133023 6 dram_wmask0[0]
port 77 nsew signal output
rlabel metal2 s 8114 132223 8170 133023 6 dram_wmask0[1]
port 78 nsew signal output
rlabel metal2 s 11150 132223 11206 133023 6 dram_wmask0[2]
port 79 nsew signal output
rlabel metal2 s 14278 132223 14334 133023 6 dram_wmask0[3]
port 80 nsew signal output
rlabel metal2 s 64602 132223 64658 133023 6 gpio_in[0]
port 81 nsew signal input
rlabel metal2 s 87878 132223 87934 133023 6 gpio_in[10]
port 82 nsew signal input
rlabel metal2 s 90178 132223 90234 133023 6 gpio_in[11]
port 83 nsew signal input
rlabel metal2 s 92478 132223 92534 133023 6 gpio_in[12]
port 84 nsew signal input
rlabel metal2 s 94870 132223 94926 133023 6 gpio_in[13]
port 85 nsew signal input
rlabel metal2 s 97170 132223 97226 133023 6 gpio_in[14]
port 86 nsew signal input
rlabel metal2 s 99470 132223 99526 133023 6 gpio_in[15]
port 87 nsew signal input
rlabel metal2 s 101862 132223 101918 133023 6 gpio_in[16]
port 88 nsew signal input
rlabel metal2 s 104162 132223 104218 133023 6 gpio_in[17]
port 89 nsew signal input
rlabel metal2 s 106462 132223 106518 133023 6 gpio_in[18]
port 90 nsew signal input
rlabel metal2 s 108762 132223 108818 133023 6 gpio_in[19]
port 91 nsew signal input
rlabel metal2 s 66994 132223 67050 133023 6 gpio_in[1]
port 92 nsew signal input
rlabel metal2 s 111154 132223 111210 133023 6 gpio_in[20]
port 93 nsew signal input
rlabel metal2 s 113454 132223 113510 133023 6 gpio_in[21]
port 94 nsew signal input
rlabel metal2 s 115754 132223 115810 133023 6 gpio_in[22]
port 95 nsew signal input
rlabel metal2 s 118054 132223 118110 133023 6 gpio_in[23]
port 96 nsew signal input
rlabel metal2 s 69294 132223 69350 133023 6 gpio_in[2]
port 97 nsew signal input
rlabel metal2 s 71594 132223 71650 133023 6 gpio_in[3]
port 98 nsew signal input
rlabel metal2 s 73894 132223 73950 133023 6 gpio_in[4]
port 99 nsew signal input
rlabel metal2 s 76286 132223 76342 133023 6 gpio_in[5]
port 100 nsew signal input
rlabel metal2 s 78586 132223 78642 133023 6 gpio_in[6]
port 101 nsew signal input
rlabel metal2 s 80886 132223 80942 133023 6 gpio_in[7]
port 102 nsew signal input
rlabel metal2 s 83186 132223 83242 133023 6 gpio_in[8]
port 103 nsew signal input
rlabel metal2 s 85578 132223 85634 133023 6 gpio_in[9]
port 104 nsew signal input
rlabel metal2 s 65430 132223 65486 133023 6 gpio_oeb[0]
port 105 nsew signal output
rlabel metal2 s 88614 132223 88670 133023 6 gpio_oeb[10]
port 106 nsew signal output
rlabel metal2 s 91006 132223 91062 133023 6 gpio_oeb[11]
port 107 nsew signal output
rlabel metal2 s 93306 132223 93362 133023 6 gpio_oeb[12]
port 108 nsew signal output
rlabel metal2 s 95606 132223 95662 133023 6 gpio_oeb[13]
port 109 nsew signal output
rlabel metal2 s 97906 132223 97962 133023 6 gpio_oeb[14]
port 110 nsew signal output
rlabel metal2 s 100298 132223 100354 133023 6 gpio_oeb[15]
port 111 nsew signal output
rlabel metal2 s 102598 132223 102654 133023 6 gpio_oeb[16]
port 112 nsew signal output
rlabel metal2 s 104898 132223 104954 133023 6 gpio_oeb[17]
port 113 nsew signal output
rlabel metal2 s 107198 132223 107254 133023 6 gpio_oeb[18]
port 114 nsew signal output
rlabel metal2 s 109590 132223 109646 133023 6 gpio_oeb[19]
port 115 nsew signal output
rlabel metal2 s 67730 132223 67786 133023 6 gpio_oeb[1]
port 116 nsew signal output
rlabel metal2 s 111890 132223 111946 133023 6 gpio_oeb[20]
port 117 nsew signal output
rlabel metal2 s 114190 132223 114246 133023 6 gpio_oeb[21]
port 118 nsew signal output
rlabel metal2 s 116582 132223 116638 133023 6 gpio_oeb[22]
port 119 nsew signal output
rlabel metal2 s 118882 132223 118938 133023 6 gpio_oeb[23]
port 120 nsew signal output
rlabel metal2 s 120446 132223 120502 133023 6 gpio_oeb[24]
port 121 nsew signal output
rlabel metal2 s 121182 132223 121238 133023 6 gpio_oeb[25]
port 122 nsew signal output
rlabel metal2 s 121918 132223 121974 133023 6 gpio_oeb[26]
port 123 nsew signal output
rlabel metal2 s 122746 132223 122802 133023 6 gpio_oeb[27]
port 124 nsew signal output
rlabel metal2 s 123482 132223 123538 133023 6 gpio_oeb[28]
port 125 nsew signal output
rlabel metal2 s 124310 132223 124366 133023 6 gpio_oeb[29]
port 126 nsew signal output
rlabel metal2 s 70030 132223 70086 133023 6 gpio_oeb[2]
port 127 nsew signal output
rlabel metal2 s 125046 132223 125102 133023 6 gpio_oeb[30]
port 128 nsew signal output
rlabel metal2 s 125874 132223 125930 133023 6 gpio_oeb[31]
port 129 nsew signal output
rlabel metal2 s 126610 132223 126666 133023 6 gpio_oeb[32]
port 130 nsew signal output
rlabel metal2 s 127346 132223 127402 133023 6 gpio_oeb[33]
port 131 nsew signal output
rlabel metal2 s 128174 132223 128230 133023 6 gpio_oeb[34]
port 132 nsew signal output
rlabel metal2 s 128910 132223 128966 133023 6 gpio_oeb[35]
port 133 nsew signal output
rlabel metal2 s 129738 132223 129794 133023 6 gpio_oeb[36]
port 134 nsew signal output
rlabel metal2 s 130474 132223 130530 133023 6 gpio_oeb[37]
port 135 nsew signal output
rlabel metal2 s 72422 132223 72478 133023 6 gpio_oeb[3]
port 136 nsew signal output
rlabel metal2 s 74722 132223 74778 133023 6 gpio_oeb[4]
port 137 nsew signal output
rlabel metal2 s 77022 132223 77078 133023 6 gpio_oeb[5]
port 138 nsew signal output
rlabel metal2 s 79322 132223 79378 133023 6 gpio_oeb[6]
port 139 nsew signal output
rlabel metal2 s 81714 132223 81770 133023 6 gpio_oeb[7]
port 140 nsew signal output
rlabel metal2 s 84014 132223 84070 133023 6 gpio_oeb[8]
port 141 nsew signal output
rlabel metal2 s 86314 132223 86370 133023 6 gpio_oeb[9]
port 142 nsew signal output
rlabel metal2 s 66166 132223 66222 133023 6 gpio_out[0]
port 143 nsew signal output
rlabel metal2 s 89442 132223 89498 133023 6 gpio_out[10]
port 144 nsew signal output
rlabel metal2 s 91742 132223 91798 133023 6 gpio_out[11]
port 145 nsew signal output
rlabel metal2 s 94042 132223 94098 133023 6 gpio_out[12]
port 146 nsew signal output
rlabel metal2 s 96434 132223 96490 133023 6 gpio_out[13]
port 147 nsew signal output
rlabel metal2 s 98734 132223 98790 133023 6 gpio_out[14]
port 148 nsew signal output
rlabel metal2 s 101034 132223 101090 133023 6 gpio_out[15]
port 149 nsew signal output
rlabel metal2 s 103334 132223 103390 133023 6 gpio_out[16]
port 150 nsew signal output
rlabel metal2 s 105726 132223 105782 133023 6 gpio_out[17]
port 151 nsew signal output
rlabel metal2 s 108026 132223 108082 133023 6 gpio_out[18]
port 152 nsew signal output
rlabel metal2 s 110326 132223 110382 133023 6 gpio_out[19]
port 153 nsew signal output
rlabel metal2 s 68466 132223 68522 133023 6 gpio_out[1]
port 154 nsew signal output
rlabel metal2 s 112626 132223 112682 133023 6 gpio_out[20]
port 155 nsew signal output
rlabel metal2 s 115018 132223 115074 133023 6 gpio_out[21]
port 156 nsew signal output
rlabel metal2 s 117318 132223 117374 133023 6 gpio_out[22]
port 157 nsew signal output
rlabel metal2 s 119618 132223 119674 133023 6 gpio_out[23]
port 158 nsew signal output
rlabel metal2 s 70858 132223 70914 133023 6 gpio_out[2]
port 159 nsew signal output
rlabel metal2 s 73158 132223 73214 133023 6 gpio_out[3]
port 160 nsew signal output
rlabel metal2 s 75458 132223 75514 133023 6 gpio_out[4]
port 161 nsew signal output
rlabel metal2 s 77850 132223 77906 133023 6 gpio_out[5]
port 162 nsew signal output
rlabel metal2 s 80150 132223 80206 133023 6 gpio_out[6]
port 163 nsew signal output
rlabel metal2 s 82450 132223 82506 133023 6 gpio_out[7]
port 164 nsew signal output
rlabel metal2 s 84750 132223 84806 133023 6 gpio_out[8]
port 165 nsew signal output
rlabel metal2 s 87142 132223 87198 133023 6 gpio_out[9]
port 166 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 iram_addr0[0]
port 167 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 iram_addr0[1]
port 168 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 iram_addr0[2]
port 169 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 iram_addr0[3]
port 170 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 iram_addr0[4]
port 171 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 iram_addr0[5]
port 172 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 iram_addr0[6]
port 173 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 iram_addr0[7]
port 174 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 iram_addr0[8]
port 175 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 iram_clk0
port 176 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 iram_csb0_A
port 177 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 iram_csb0_B
port 178 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 iram_din0[0]
port 179 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 iram_din0[10]
port 180 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 iram_din0[11]
port 181 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 iram_din0[12]
port 182 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 iram_din0[13]
port 183 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 iram_din0[14]
port 184 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 iram_din0[15]
port 185 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 iram_din0[16]
port 186 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 iram_din0[17]
port 187 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 iram_din0[18]
port 188 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 iram_din0[19]
port 189 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 iram_din0[1]
port 190 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 iram_din0[20]
port 191 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 iram_din0[21]
port 192 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 iram_din0[22]
port 193 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 iram_din0[23]
port 194 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 iram_din0[24]
port 195 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 iram_din0[25]
port 196 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 iram_din0[26]
port 197 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 iram_din0[27]
port 198 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 iram_din0[28]
port 199 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 iram_din0[29]
port 200 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 iram_din0[2]
port 201 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 iram_din0[30]
port 202 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 iram_din0[31]
port 203 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 iram_din0[3]
port 204 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 iram_din0[4]
port 205 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 iram_din0[5]
port 206 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 iram_din0[6]
port 207 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 iram_din0[7]
port 208 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 iram_din0[8]
port 209 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 iram_din0[9]
port 210 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 iram_dout0_A[0]
port 211 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 iram_dout0_A[10]
port 212 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 iram_dout0_A[11]
port 213 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 iram_dout0_A[12]
port 214 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 iram_dout0_A[13]
port 215 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 iram_dout0_A[14]
port 216 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 iram_dout0_A[15]
port 217 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 iram_dout0_A[16]
port 218 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 iram_dout0_A[17]
port 219 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 iram_dout0_A[18]
port 220 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 iram_dout0_A[19]
port 221 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 iram_dout0_A[1]
port 222 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 iram_dout0_A[20]
port 223 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 iram_dout0_A[21]
port 224 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 iram_dout0_A[22]
port 225 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 iram_dout0_A[23]
port 226 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 iram_dout0_A[24]
port 227 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 iram_dout0_A[25]
port 228 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 iram_dout0_A[26]
port 229 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 iram_dout0_A[27]
port 230 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 iram_dout0_A[28]
port 231 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 iram_dout0_A[29]
port 232 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 iram_dout0_A[2]
port 233 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 iram_dout0_A[30]
port 234 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 iram_dout0_A[31]
port 235 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 iram_dout0_A[3]
port 236 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 iram_dout0_A[4]
port 237 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 iram_dout0_A[5]
port 238 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 iram_dout0_A[6]
port 239 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 iram_dout0_A[7]
port 240 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 iram_dout0_A[8]
port 241 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 iram_dout0_A[9]
port 242 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 iram_dout0_B[0]
port 243 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 iram_dout0_B[10]
port 244 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 iram_dout0_B[11]
port 245 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 iram_dout0_B[12]
port 246 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 iram_dout0_B[13]
port 247 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 iram_dout0_B[14]
port 248 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 iram_dout0_B[15]
port 249 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 iram_dout0_B[16]
port 250 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 iram_dout0_B[17]
port 251 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 iram_dout0_B[18]
port 252 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 iram_dout0_B[19]
port 253 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 iram_dout0_B[1]
port 254 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 iram_dout0_B[20]
port 255 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 iram_dout0_B[21]
port 256 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 iram_dout0_B[22]
port 257 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 iram_dout0_B[23]
port 258 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 iram_dout0_B[24]
port 259 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 iram_dout0_B[25]
port 260 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 iram_dout0_B[26]
port 261 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 iram_dout0_B[27]
port 262 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 iram_dout0_B[28]
port 263 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 iram_dout0_B[29]
port 264 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 iram_dout0_B[2]
port 265 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 iram_dout0_B[30]
port 266 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 iram_dout0_B[31]
port 267 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 iram_dout0_B[3]
port 268 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 iram_dout0_B[4]
port 269 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 iram_dout0_B[5]
port 270 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 iram_dout0_B[6]
port 271 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 iram_dout0_B[7]
port 272 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 iram_dout0_B[8]
port 273 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 iram_dout0_B[9]
port 274 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 iram_web0
port 275 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 iram_wmask0[0]
port 276 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 iram_wmask0[1]
port 277 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 iram_wmask0[2]
port 278 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 iram_wmask0[3]
port 279 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 la_data_in[0]
port 280 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[100]
port 281 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[101]
port 282 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[102]
port 283 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[103]
port 284 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[104]
port 285 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[105]
port 286 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[106]
port 287 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_data_in[107]
port 288 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[108]
port 289 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[109]
port 290 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[10]
port 291 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[110]
port 292 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[111]
port 293 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[112]
port 294 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[113]
port 295 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_data_in[114]
port 296 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[115]
port 297 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[116]
port 298 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[117]
port 299 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[118]
port 300 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[119]
port 301 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[11]
port 302 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[120]
port 303 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[121]
port 304 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_data_in[122]
port 305 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[123]
port 306 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[124]
port 307 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[125]
port 308 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[126]
port 309 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[127]
port 310 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[12]
port 311 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[13]
port 312 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_data_in[14]
port 313 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[15]
port 314 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in[16]
port 315 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[17]
port 316 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_in[18]
port 317 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[19]
port 318 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_data_in[1]
port 319 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[20]
port 320 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[21]
port 321 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_data_in[22]
port 322 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[23]
port 323 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_in[24]
port 324 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_in[25]
port 325 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[26]
port 326 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[27]
port 327 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[28]
port 328 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[29]
port 329 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_data_in[2]
port 330 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[30]
port 331 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[31]
port 332 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[32]
port 333 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[33]
port 334 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[34]
port 335 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[35]
port 336 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[36]
port 337 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[37]
port 338 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[38]
port 339 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[39]
port 340 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_data_in[3]
port 341 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_data_in[40]
port 342 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[41]
port 343 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[42]
port 344 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[43]
port 345 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in[44]
port 346 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[45]
port 347 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[46]
port 348 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[47]
port 349 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[48]
port 350 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[49]
port 351 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[4]
port 352 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[50]
port 353 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[51]
port 354 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[52]
port 355 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[53]
port 356 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[54]
port 357 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[55]
port 358 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_data_in[56]
port 359 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[57]
port 360 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[58]
port 361 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[59]
port 362 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_data_in[5]
port 363 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[60]
port 364 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[61]
port 365 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[62]
port 366 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[63]
port 367 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[64]
port 368 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[65]
port 369 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_data_in[66]
port 370 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[67]
port 371 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[68]
port 372 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[69]
port 373 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[6]
port 374 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[70]
port 375 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[71]
port 376 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[72]
port 377 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[73]
port 378 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[74]
port 379 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[75]
port 380 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[76]
port 381 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_data_in[77]
port 382 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[78]
port 383 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[79]
port 384 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[7]
port 385 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_data_in[80]
port 386 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[81]
port 387 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[82]
port 388 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[83]
port 389 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[84]
port 390 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[85]
port 391 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[86]
port 392 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[87]
port 393 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_data_in[88]
port 394 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[89]
port 395 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_data_in[8]
port 396 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[90]
port 397 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_data_in[91]
port 398 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[92]
port 399 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[93]
port 400 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[94]
port 401 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[95]
port 402 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[96]
port 403 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[97]
port 404 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[98]
port 405 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[99]
port 406 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[9]
port 407 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_data_out[0]
port 408 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[100]
port 409 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 la_data_out[101]
port 410 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[102]
port 411 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[103]
port 412 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[104]
port 413 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[105]
port 414 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[106]
port 415 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[107]
port 416 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[108]
port 417 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[109]
port 418 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 la_data_out[10]
port 419 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[110]
port 420 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[111]
port 421 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[112]
port 422 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[113]
port 423 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 la_data_out[114]
port 424 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[115]
port 425 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[116]
port 426 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[117]
port 427 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[118]
port 428 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 la_data_out[119]
port 429 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 la_data_out[11]
port 430 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 la_data_out[120]
port 431 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[121]
port 432 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[122]
port 433 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[123]
port 434 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 la_data_out[124]
port 435 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[125]
port 436 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[126]
port 437 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 la_data_out[127]
port 438 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 la_data_out[12]
port 439 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 la_data_out[13]
port 440 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 la_data_out[14]
port 441 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[15]
port 442 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 la_data_out[16]
port 443 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 la_data_out[17]
port 444 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 la_data_out[18]
port 445 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 la_data_out[19]
port 446 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 la_data_out[1]
port 447 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[20]
port 448 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 la_data_out[21]
port 449 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[22]
port 450 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[23]
port 451 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[24]
port 452 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 la_data_out[25]
port 453 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[26]
port 454 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[27]
port 455 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[28]
port 456 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[29]
port 457 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 la_data_out[2]
port 458 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[30]
port 459 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 la_data_out[31]
port 460 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_data_out[32]
port 461 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[33]
port 462 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[34]
port 463 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[35]
port 464 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 la_data_out[36]
port 465 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[37]
port 466 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[38]
port 467 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[39]
port 468 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 la_data_out[3]
port 469 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[40]
port 470 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[41]
port 471 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[42]
port 472 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[43]
port 473 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[44]
port 474 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[45]
port 475 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[46]
port 476 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[47]
port 477 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[48]
port 478 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[49]
port 479 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 la_data_out[4]
port 480 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[50]
port 481 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 la_data_out[51]
port 482 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[52]
port 483 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[53]
port 484 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[54]
port 485 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[55]
port 486 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[56]
port 487 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[57]
port 488 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[58]
port 489 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[59]
port 490 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 la_data_out[5]
port 491 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[60]
port 492 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[61]
port 493 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[62]
port 494 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[63]
port 495 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[64]
port 496 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[65]
port 497 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[66]
port 498 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[67]
port 499 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 la_data_out[68]
port 500 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[69]
port 501 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 la_data_out[6]
port 502 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[70]
port 503 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[71]
port 504 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[72]
port 505 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[73]
port 506 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[74]
port 507 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[75]
port 508 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[76]
port 509 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[77]
port 510 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[78]
port 511 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[79]
port 512 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 la_data_out[7]
port 513 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[80]
port 514 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 la_data_out[81]
port 515 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[82]
port 516 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[83]
port 517 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[84]
port 518 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[85]
port 519 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 la_data_out[86]
port 520 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[87]
port 521 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[88]
port 522 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[89]
port 523 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 la_data_out[8]
port 524 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 la_data_out[90]
port 525 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 la_data_out[91]
port 526 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[92]
port 527 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[93]
port 528 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[94]
port 529 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[95]
port 530 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 la_data_out[96]
port 531 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[97]
port 532 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[98]
port 533 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[99]
port 534 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[9]
port 535 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 la_oenb[0]
port 536 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[100]
port 537 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[101]
port 538 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[102]
port 539 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[103]
port 540 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[104]
port 541 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[105]
port 542 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[106]
port 543 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[107]
port 544 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[108]
port 545 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_oenb[109]
port 546 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_oenb[10]
port 547 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[110]
port 548 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[111]
port 549 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[112]
port 550 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[113]
port 551 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oenb[114]
port 552 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_oenb[115]
port 553 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[116]
port 554 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[117]
port 555 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[118]
port 556 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_oenb[119]
port 557 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_oenb[11]
port 558 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[120]
port 559 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_oenb[121]
port 560 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_oenb[122]
port 561 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_oenb[123]
port 562 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oenb[124]
port 563 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_oenb[125]
port 564 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_oenb[126]
port 565 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[127]
port 566 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_oenb[12]
port 567 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_oenb[13]
port 568 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_oenb[14]
port 569 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[15]
port 570 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_oenb[16]
port 571 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_oenb[17]
port 572 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[18]
port 573 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[19]
port 574 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 la_oenb[1]
port 575 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[20]
port 576 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_oenb[21]
port 577 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[22]
port 578 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[23]
port 579 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[24]
port 580 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_oenb[25]
port 581 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[26]
port 582 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[27]
port 583 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_oenb[28]
port 584 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[29]
port 585 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_oenb[2]
port 586 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[30]
port 587 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[31]
port 588 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[32]
port 589 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[33]
port 590 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_oenb[34]
port 591 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[35]
port 592 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_oenb[36]
port 593 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[37]
port 594 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[38]
port 595 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[39]
port 596 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[3]
port 597 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[40]
port 598 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[41]
port 599 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[42]
port 600 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_oenb[43]
port 601 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[44]
port 602 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[45]
port 603 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_oenb[46]
port 604 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[47]
port 605 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[48]
port 606 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_oenb[49]
port 607 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_oenb[4]
port 608 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[50]
port 609 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[51]
port 610 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[52]
port 611 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[53]
port 612 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oenb[54]
port 613 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[55]
port 614 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[56]
port 615 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[57]
port 616 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[58]
port 617 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[59]
port 618 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_oenb[5]
port 619 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_oenb[60]
port 620 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[61]
port 621 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[62]
port 622 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_oenb[63]
port 623 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_oenb[64]
port 624 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[65]
port 625 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[66]
port 626 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[67]
port 627 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oenb[68]
port 628 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_oenb[69]
port 629 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_oenb[6]
port 630 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oenb[70]
port 631 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_oenb[71]
port 632 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[72]
port 633 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_oenb[73]
port 634 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[74]
port 635 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[75]
port 636 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[76]
port 637 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[77]
port 638 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[78]
port 639 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[79]
port 640 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[7]
port 641 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[80]
port 642 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[81]
port 643 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[82]
port 644 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[83]
port 645 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[84]
port 646 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[85]
port 647 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_oenb[86]
port 648 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[87]
port 649 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[88]
port 650 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[89]
port 651 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[8]
port 652 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[90]
port 653 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[91]
port 654 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[92]
port 655 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[93]
port 656 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[94]
port 657 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[95]
port 658 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[96]
port 659 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[97]
port 660 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[98]
port 661 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[99]
port 662 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[9]
port 663 nsew signal input
rlabel metal2 s 62302 132223 62358 133023 6 user_irq[0]
port 664 nsew signal output
rlabel metal2 s 63130 132223 63186 133023 6 user_irq[1]
port 665 nsew signal output
rlabel metal2 s 63866 132223 63922 133023 6 user_irq[2]
port 666 nsew signal output
rlabel metal4 s 4208 2128 4528 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 669 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 670 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 671 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[0]
port 672 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[10]
port 673 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[11]
port 674 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[12]
port 675 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_adr_i[13]
port 676 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[14]
port 677 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[15]
port 678 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[16]
port 679 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[17]
port 680 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[18]
port 681 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[19]
port 682 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[1]
port 683 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_adr_i[20]
port 684 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[21]
port 685 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[22]
port 686 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[23]
port 687 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[24]
port 688 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[25]
port 689 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[26]
port 690 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[27]
port 691 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[28]
port 692 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[29]
port 693 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_adr_i[2]
port 694 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[30]
port 695 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[31]
port 696 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[3]
port 697 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[4]
port 698 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[5]
port 699 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[6]
port 700 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[7]
port 701 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[8]
port 702 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[9]
port 703 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 704 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_i[0]
port 705 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[10]
port 706 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[11]
port 707 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[12]
port 708 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[13]
port 709 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[14]
port 710 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[15]
port 711 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[16]
port 712 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_i[17]
port 713 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_i[18]
port 714 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[19]
port 715 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_i[1]
port 716 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_i[20]
port 717 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[21]
port 718 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[22]
port 719 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[23]
port 720 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[24]
port 721 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[25]
port 722 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[26]
port 723 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_i[27]
port 724 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_i[28]
port 725 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[29]
port 726 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[2]
port 727 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[30]
port 728 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[31]
port 729 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[3]
port 730 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_i[4]
port 731 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[5]
port 732 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[6]
port 733 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[7]
port 734 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[8]
port 735 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[9]
port 736 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_o[0]
port 737 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[10]
port 738 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[11]
port 739 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[12]
port 740 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[13]
port 741 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[14]
port 742 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[15]
port 743 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[16]
port 744 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[17]
port 745 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[18]
port 746 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_o[19]
port 747 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[1]
port 748 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_o[20]
port 749 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_o[21]
port 750 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[22]
port 751 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[23]
port 752 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[24]
port 753 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[25]
port 754 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[26]
port 755 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[27]
port 756 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[28]
port 757 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[29]
port 758 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_o[2]
port 759 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[30]
port 760 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[31]
port 761 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[3]
port 762 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_o[4]
port 763 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[5]
port 764 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[6]
port 765 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[7]
port 766 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[8]
port 767 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[9]
port 768 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 wbs_sel_i[0]
port 769 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_sel_i[1]
port 770 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[2]
port 771 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_sel_i[3]
port 772 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_stb_i
port 773 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 774 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 130879 133023
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 43975250
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc/openlane/rvj1_caravel_soc/runs/rvj1_caravel_soc/results/signoff/rvj1_caravel_soc.magic.gds
string GDS_START 1228438
<< end >>

