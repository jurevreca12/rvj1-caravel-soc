magic
tech sky130A
magscale 1 2
timestamp 1653847779
<< obsli1 >>
rect 1104 2159 118588 119697
<< obsm1 >>
rect 106 416 119678 119808
<< metal2 >>
rect 294 121102 350 121902
rect 846 121102 902 121902
rect 1490 121102 1546 121902
rect 2042 121102 2098 121902
rect 2686 121102 2742 121902
rect 3330 121102 3386 121902
rect 3882 121102 3938 121902
rect 4526 121102 4582 121902
rect 5078 121102 5134 121902
rect 5722 121102 5778 121902
rect 6366 121102 6422 121902
rect 6918 121102 6974 121902
rect 7562 121102 7618 121902
rect 8114 121102 8170 121902
rect 8758 121102 8814 121902
rect 9402 121102 9458 121902
rect 9954 121102 10010 121902
rect 10598 121102 10654 121902
rect 11150 121102 11206 121902
rect 11794 121102 11850 121902
rect 12438 121102 12494 121902
rect 12990 121102 13046 121902
rect 13634 121102 13690 121902
rect 14278 121102 14334 121902
rect 14830 121102 14886 121902
rect 15474 121102 15530 121902
rect 16026 121102 16082 121902
rect 16670 121102 16726 121902
rect 17314 121102 17370 121902
rect 17866 121102 17922 121902
rect 18510 121102 18566 121902
rect 19062 121102 19118 121902
rect 19706 121102 19762 121902
rect 20350 121102 20406 121902
rect 20902 121102 20958 121902
rect 21546 121102 21602 121902
rect 22098 121102 22154 121902
rect 22742 121102 22798 121902
rect 23386 121102 23442 121902
rect 23938 121102 23994 121902
rect 24582 121102 24638 121902
rect 25134 121102 25190 121902
rect 25778 121102 25834 121902
rect 26422 121102 26478 121902
rect 26974 121102 27030 121902
rect 27618 121102 27674 121902
rect 28262 121102 28318 121902
rect 28814 121102 28870 121902
rect 29458 121102 29514 121902
rect 30010 121102 30066 121902
rect 30654 121102 30710 121902
rect 31298 121102 31354 121902
rect 31850 121102 31906 121902
rect 32494 121102 32550 121902
rect 33046 121102 33102 121902
rect 33690 121102 33746 121902
rect 34334 121102 34390 121902
rect 34886 121102 34942 121902
rect 35530 121102 35586 121902
rect 36082 121102 36138 121902
rect 36726 121102 36782 121902
rect 37370 121102 37426 121902
rect 37922 121102 37978 121902
rect 38566 121102 38622 121902
rect 39118 121102 39174 121902
rect 39762 121102 39818 121902
rect 40406 121102 40462 121902
rect 40958 121102 41014 121902
rect 41602 121102 41658 121902
rect 42246 121102 42302 121902
rect 42798 121102 42854 121902
rect 43442 121102 43498 121902
rect 43994 121102 44050 121902
rect 44638 121102 44694 121902
rect 45282 121102 45338 121902
rect 45834 121102 45890 121902
rect 46478 121102 46534 121902
rect 47030 121102 47086 121902
rect 47674 121102 47730 121902
rect 48318 121102 48374 121902
rect 48870 121102 48926 121902
rect 49514 121102 49570 121902
rect 50066 121102 50122 121902
rect 50710 121102 50766 121902
rect 51354 121102 51410 121902
rect 51906 121102 51962 121902
rect 52550 121102 52606 121902
rect 53102 121102 53158 121902
rect 53746 121102 53802 121902
rect 54390 121102 54446 121902
rect 54942 121102 54998 121902
rect 55586 121102 55642 121902
rect 56230 121102 56286 121902
rect 56782 121102 56838 121902
rect 57426 121102 57482 121902
rect 57978 121102 58034 121902
rect 58622 121102 58678 121902
rect 59266 121102 59322 121902
rect 59818 121102 59874 121902
rect 60462 121102 60518 121902
rect 61014 121102 61070 121902
rect 61658 121102 61714 121902
rect 62302 121102 62358 121902
rect 62854 121102 62910 121902
rect 63498 121102 63554 121902
rect 64050 121102 64106 121902
rect 64694 121102 64750 121902
rect 65338 121102 65394 121902
rect 65890 121102 65946 121902
rect 66534 121102 66590 121902
rect 67178 121102 67234 121902
rect 67730 121102 67786 121902
rect 68374 121102 68430 121902
rect 68926 121102 68982 121902
rect 69570 121102 69626 121902
rect 70214 121102 70270 121902
rect 70766 121102 70822 121902
rect 71410 121102 71466 121902
rect 71962 121102 72018 121902
rect 72606 121102 72662 121902
rect 73250 121102 73306 121902
rect 73802 121102 73858 121902
rect 74446 121102 74502 121902
rect 74998 121102 75054 121902
rect 75642 121102 75698 121902
rect 76286 121102 76342 121902
rect 76838 121102 76894 121902
rect 77482 121102 77538 121902
rect 78034 121102 78090 121902
rect 78678 121102 78734 121902
rect 79322 121102 79378 121902
rect 79874 121102 79930 121902
rect 80518 121102 80574 121902
rect 81162 121102 81218 121902
rect 81714 121102 81770 121902
rect 82358 121102 82414 121902
rect 82910 121102 82966 121902
rect 83554 121102 83610 121902
rect 84198 121102 84254 121902
rect 84750 121102 84806 121902
rect 85394 121102 85450 121902
rect 85946 121102 86002 121902
rect 86590 121102 86646 121902
rect 87234 121102 87290 121902
rect 87786 121102 87842 121902
rect 88430 121102 88486 121902
rect 88982 121102 89038 121902
rect 89626 121102 89682 121902
rect 90270 121102 90326 121902
rect 90822 121102 90878 121902
rect 91466 121102 91522 121902
rect 92018 121102 92074 121902
rect 92662 121102 92718 121902
rect 93306 121102 93362 121902
rect 93858 121102 93914 121902
rect 94502 121102 94558 121902
rect 95146 121102 95202 121902
rect 95698 121102 95754 121902
rect 96342 121102 96398 121902
rect 96894 121102 96950 121902
rect 97538 121102 97594 121902
rect 98182 121102 98238 121902
rect 98734 121102 98790 121902
rect 99378 121102 99434 121902
rect 99930 121102 99986 121902
rect 100574 121102 100630 121902
rect 101218 121102 101274 121902
rect 101770 121102 101826 121902
rect 102414 121102 102470 121902
rect 102966 121102 103022 121902
rect 103610 121102 103666 121902
rect 104254 121102 104310 121902
rect 104806 121102 104862 121902
rect 105450 121102 105506 121902
rect 106002 121102 106058 121902
rect 106646 121102 106702 121902
rect 107290 121102 107346 121902
rect 107842 121102 107898 121902
rect 108486 121102 108542 121902
rect 109130 121102 109186 121902
rect 109682 121102 109738 121902
rect 110326 121102 110382 121902
rect 110878 121102 110934 121902
rect 111522 121102 111578 121902
rect 112166 121102 112222 121902
rect 112718 121102 112774 121902
rect 113362 121102 113418 121902
rect 113914 121102 113970 121902
rect 114558 121102 114614 121902
rect 115202 121102 115258 121902
rect 115754 121102 115810 121902
rect 116398 121102 116454 121902
rect 116950 121102 117006 121902
rect 117594 121102 117650 121902
rect 118238 121102 118294 121902
rect 118790 121102 118846 121902
rect 119434 121102 119490 121902
rect 18 0 74 800
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5262 0 5318 800
rect 5446 0 5502 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 18050 0 18106 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46754 0 46810 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66074 0 66130 800
rect 66258 0 66314 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67086 0 67142 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74354 0 74410 800
rect 74538 0 74594 800
rect 74722 0 74778 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75826 0 75882 800
rect 76010 0 76066 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79690 0 79746 800
rect 79874 0 79930 800
rect 80058 0 80114 800
rect 80242 0 80298 800
rect 80426 0 80482 800
rect 80610 0 80666 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 83922 0 83978 800
rect 84106 0 84162 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85578 0 85634 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86130 0 86186 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86774 0 86830 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89258 0 89314 800
rect 89442 0 89498 800
rect 89626 0 89682 800
rect 89810 0 89866 800
rect 89994 0 90050 800
rect 90178 0 90234 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91006 0 91062 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92478 0 92534 800
rect 92662 0 92718 800
rect 92846 0 92902 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93490 0 93546 800
rect 93674 0 93730 800
rect 93858 0 93914 800
rect 94042 0 94098 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95146 0 95202 800
rect 95330 0 95386 800
rect 95514 0 95570 800
rect 95698 0 95754 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96158 0 96214 800
rect 96342 0 96398 800
rect 96526 0 96582 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97078 0 97134 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98182 0 98238 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99194 0 99250 800
rect 99378 0 99434 800
rect 99562 0 99618 800
rect 99746 0 99802 800
rect 99930 0 99986 800
rect 100114 0 100170 800
rect 100298 0 100354 800
rect 100482 0 100538 800
rect 100574 0 100630 800
rect 100758 0 100814 800
rect 100942 0 100998 800
rect 101126 0 101182 800
rect 101310 0 101366 800
rect 101494 0 101550 800
rect 101678 0 101734 800
rect 101862 0 101918 800
rect 102046 0 102102 800
rect 102230 0 102286 800
rect 102414 0 102470 800
rect 102598 0 102654 800
rect 102782 0 102838 800
rect 102966 0 103022 800
rect 103058 0 103114 800
rect 103242 0 103298 800
rect 103426 0 103482 800
rect 103610 0 103666 800
rect 103794 0 103850 800
rect 103978 0 104034 800
rect 104162 0 104218 800
rect 104346 0 104402 800
rect 104530 0 104586 800
rect 104714 0 104770 800
rect 104898 0 104954 800
rect 105082 0 105138 800
rect 105266 0 105322 800
rect 105358 0 105414 800
rect 105542 0 105598 800
rect 105726 0 105782 800
rect 105910 0 105966 800
rect 106094 0 106150 800
rect 106278 0 106334 800
rect 106462 0 106518 800
rect 106646 0 106702 800
rect 106830 0 106886 800
rect 107014 0 107070 800
rect 107198 0 107254 800
rect 107382 0 107438 800
rect 107566 0 107622 800
rect 107750 0 107806 800
rect 107842 0 107898 800
rect 108026 0 108082 800
rect 108210 0 108266 800
rect 108394 0 108450 800
rect 108578 0 108634 800
rect 108762 0 108818 800
rect 108946 0 109002 800
rect 109130 0 109186 800
rect 109314 0 109370 800
rect 109498 0 109554 800
rect 109682 0 109738 800
rect 109866 0 109922 800
rect 110050 0 110106 800
rect 110142 0 110198 800
rect 110326 0 110382 800
rect 110510 0 110566 800
rect 110694 0 110750 800
rect 110878 0 110934 800
rect 111062 0 111118 800
rect 111246 0 111302 800
rect 111430 0 111486 800
rect 111614 0 111670 800
rect 111798 0 111854 800
rect 111982 0 112038 800
rect 112166 0 112222 800
rect 112350 0 112406 800
rect 112534 0 112590 800
rect 112626 0 112682 800
rect 112810 0 112866 800
rect 112994 0 113050 800
rect 113178 0 113234 800
rect 113362 0 113418 800
rect 113546 0 113602 800
rect 113730 0 113786 800
rect 113914 0 113970 800
rect 114098 0 114154 800
rect 114282 0 114338 800
rect 114466 0 114522 800
rect 114650 0 114706 800
rect 114834 0 114890 800
rect 114926 0 114982 800
rect 115110 0 115166 800
rect 115294 0 115350 800
rect 115478 0 115534 800
rect 115662 0 115718 800
rect 115846 0 115902 800
rect 116030 0 116086 800
rect 116214 0 116270 800
rect 116398 0 116454 800
rect 116582 0 116638 800
rect 116766 0 116822 800
rect 116950 0 117006 800
rect 117134 0 117190 800
rect 117318 0 117374 800
rect 117410 0 117466 800
rect 117594 0 117650 800
rect 117778 0 117834 800
rect 117962 0 118018 800
rect 118146 0 118202 800
rect 118330 0 118386 800
rect 118514 0 118570 800
rect 118698 0 118754 800
rect 118882 0 118938 800
rect 119066 0 119122 800
rect 119250 0 119306 800
rect 119434 0 119490 800
rect 119618 0 119674 800
<< obsm2 >>
rect 18 121046 238 121258
rect 406 121046 790 121258
rect 958 121046 1434 121258
rect 1602 121046 1986 121258
rect 2154 121046 2630 121258
rect 2798 121046 3274 121258
rect 3442 121046 3826 121258
rect 3994 121046 4470 121258
rect 4638 121046 5022 121258
rect 5190 121046 5666 121258
rect 5834 121046 6310 121258
rect 6478 121046 6862 121258
rect 7030 121046 7506 121258
rect 7674 121046 8058 121258
rect 8226 121046 8702 121258
rect 8870 121046 9346 121258
rect 9514 121046 9898 121258
rect 10066 121046 10542 121258
rect 10710 121046 11094 121258
rect 11262 121046 11738 121258
rect 11906 121046 12382 121258
rect 12550 121046 12934 121258
rect 13102 121046 13578 121258
rect 13746 121046 14222 121258
rect 14390 121046 14774 121258
rect 14942 121046 15418 121258
rect 15586 121046 15970 121258
rect 16138 121046 16614 121258
rect 16782 121046 17258 121258
rect 17426 121046 17810 121258
rect 17978 121046 18454 121258
rect 18622 121046 19006 121258
rect 19174 121046 19650 121258
rect 19818 121046 20294 121258
rect 20462 121046 20846 121258
rect 21014 121046 21490 121258
rect 21658 121046 22042 121258
rect 22210 121046 22686 121258
rect 22854 121046 23330 121258
rect 23498 121046 23882 121258
rect 24050 121046 24526 121258
rect 24694 121046 25078 121258
rect 25246 121046 25722 121258
rect 25890 121046 26366 121258
rect 26534 121046 26918 121258
rect 27086 121046 27562 121258
rect 27730 121046 28206 121258
rect 28374 121046 28758 121258
rect 28926 121046 29402 121258
rect 29570 121046 29954 121258
rect 30122 121046 30598 121258
rect 30766 121046 31242 121258
rect 31410 121046 31794 121258
rect 31962 121046 32438 121258
rect 32606 121046 32990 121258
rect 33158 121046 33634 121258
rect 33802 121046 34278 121258
rect 34446 121046 34830 121258
rect 34998 121046 35474 121258
rect 35642 121046 36026 121258
rect 36194 121046 36670 121258
rect 36838 121046 37314 121258
rect 37482 121046 37866 121258
rect 38034 121046 38510 121258
rect 38678 121046 39062 121258
rect 39230 121046 39706 121258
rect 39874 121046 40350 121258
rect 40518 121046 40902 121258
rect 41070 121046 41546 121258
rect 41714 121046 42190 121258
rect 42358 121046 42742 121258
rect 42910 121046 43386 121258
rect 43554 121046 43938 121258
rect 44106 121046 44582 121258
rect 44750 121046 45226 121258
rect 45394 121046 45778 121258
rect 45946 121046 46422 121258
rect 46590 121046 46974 121258
rect 47142 121046 47618 121258
rect 47786 121046 48262 121258
rect 48430 121046 48814 121258
rect 48982 121046 49458 121258
rect 49626 121046 50010 121258
rect 50178 121046 50654 121258
rect 50822 121046 51298 121258
rect 51466 121046 51850 121258
rect 52018 121046 52494 121258
rect 52662 121046 53046 121258
rect 53214 121046 53690 121258
rect 53858 121046 54334 121258
rect 54502 121046 54886 121258
rect 55054 121046 55530 121258
rect 55698 121046 56174 121258
rect 56342 121046 56726 121258
rect 56894 121046 57370 121258
rect 57538 121046 57922 121258
rect 58090 121046 58566 121258
rect 58734 121046 59210 121258
rect 59378 121046 59762 121258
rect 59930 121046 60406 121258
rect 60574 121046 60958 121258
rect 61126 121046 61602 121258
rect 61770 121046 62246 121258
rect 62414 121046 62798 121258
rect 62966 121046 63442 121258
rect 63610 121046 63994 121258
rect 64162 121046 64638 121258
rect 64806 121046 65282 121258
rect 65450 121046 65834 121258
rect 66002 121046 66478 121258
rect 66646 121046 67122 121258
rect 67290 121046 67674 121258
rect 67842 121046 68318 121258
rect 68486 121046 68870 121258
rect 69038 121046 69514 121258
rect 69682 121046 70158 121258
rect 70326 121046 70710 121258
rect 70878 121046 71354 121258
rect 71522 121046 71906 121258
rect 72074 121046 72550 121258
rect 72718 121046 73194 121258
rect 73362 121046 73746 121258
rect 73914 121046 74390 121258
rect 74558 121046 74942 121258
rect 75110 121046 75586 121258
rect 75754 121046 76230 121258
rect 76398 121046 76782 121258
rect 76950 121046 77426 121258
rect 77594 121046 77978 121258
rect 78146 121046 78622 121258
rect 78790 121046 79266 121258
rect 79434 121046 79818 121258
rect 79986 121046 80462 121258
rect 80630 121046 81106 121258
rect 81274 121046 81658 121258
rect 81826 121046 82302 121258
rect 82470 121046 82854 121258
rect 83022 121046 83498 121258
rect 83666 121046 84142 121258
rect 84310 121046 84694 121258
rect 84862 121046 85338 121258
rect 85506 121046 85890 121258
rect 86058 121046 86534 121258
rect 86702 121046 87178 121258
rect 87346 121046 87730 121258
rect 87898 121046 88374 121258
rect 88542 121046 88926 121258
rect 89094 121046 89570 121258
rect 89738 121046 90214 121258
rect 90382 121046 90766 121258
rect 90934 121046 91410 121258
rect 91578 121046 91962 121258
rect 92130 121046 92606 121258
rect 92774 121046 93250 121258
rect 93418 121046 93802 121258
rect 93970 121046 94446 121258
rect 94614 121046 95090 121258
rect 95258 121046 95642 121258
rect 95810 121046 96286 121258
rect 96454 121046 96838 121258
rect 97006 121046 97482 121258
rect 97650 121046 98126 121258
rect 98294 121046 98678 121258
rect 98846 121046 99322 121258
rect 99490 121046 99874 121258
rect 100042 121046 100518 121258
rect 100686 121046 101162 121258
rect 101330 121046 101714 121258
rect 101882 121046 102358 121258
rect 102526 121046 102910 121258
rect 103078 121046 103554 121258
rect 103722 121046 104198 121258
rect 104366 121046 104750 121258
rect 104918 121046 105394 121258
rect 105562 121046 105946 121258
rect 106114 121046 106590 121258
rect 106758 121046 107234 121258
rect 107402 121046 107786 121258
rect 107954 121046 108430 121258
rect 108598 121046 109074 121258
rect 109242 121046 109626 121258
rect 109794 121046 110270 121258
rect 110438 121046 110822 121258
rect 110990 121046 111466 121258
rect 111634 121046 112110 121258
rect 112278 121046 112662 121258
rect 112830 121046 113306 121258
rect 113474 121046 113858 121258
rect 114026 121046 114502 121258
rect 114670 121046 115146 121258
rect 115314 121046 115698 121258
rect 115866 121046 116342 121258
rect 116510 121046 116894 121258
rect 117062 121046 117538 121258
rect 117706 121046 118182 121258
rect 118350 121046 118734 121258
rect 118902 121046 119378 121258
rect 119546 121046 119672 121258
rect 18 856 119672 121046
rect 222 303 238 856
rect 406 303 422 856
rect 590 303 606 856
rect 774 303 790 856
rect 958 303 974 856
rect 1142 303 1158 856
rect 1326 303 1342 856
rect 1510 303 1526 856
rect 1694 303 1710 856
rect 1878 303 1894 856
rect 2062 303 2078 856
rect 2246 303 2262 856
rect 2522 303 2538 856
rect 2706 303 2722 856
rect 2890 303 2906 856
rect 3074 303 3090 856
rect 3258 303 3274 856
rect 3442 303 3458 856
rect 3626 303 3642 856
rect 3810 303 3826 856
rect 3994 303 4010 856
rect 4178 303 4194 856
rect 4362 303 4378 856
rect 4546 303 4562 856
rect 4730 303 4746 856
rect 5006 303 5022 856
rect 5190 303 5206 856
rect 5374 303 5390 856
rect 5558 303 5574 856
rect 5742 303 5758 856
rect 5926 303 5942 856
rect 6110 303 6126 856
rect 6294 303 6310 856
rect 6478 303 6494 856
rect 6662 303 6678 856
rect 6846 303 6862 856
rect 7030 303 7046 856
rect 7306 303 7322 856
rect 7490 303 7506 856
rect 7674 303 7690 856
rect 7858 303 7874 856
rect 8042 303 8058 856
rect 8226 303 8242 856
rect 8410 303 8426 856
rect 8594 303 8610 856
rect 8778 303 8794 856
rect 8962 303 8978 856
rect 9146 303 9162 856
rect 9330 303 9346 856
rect 9514 303 9530 856
rect 9790 303 9806 856
rect 9974 303 9990 856
rect 10158 303 10174 856
rect 10342 303 10358 856
rect 10526 303 10542 856
rect 10710 303 10726 856
rect 10894 303 10910 856
rect 11078 303 11094 856
rect 11262 303 11278 856
rect 11446 303 11462 856
rect 11630 303 11646 856
rect 11814 303 11830 856
rect 12090 303 12106 856
rect 12274 303 12290 856
rect 12458 303 12474 856
rect 12642 303 12658 856
rect 12826 303 12842 856
rect 13010 303 13026 856
rect 13194 303 13210 856
rect 13378 303 13394 856
rect 13562 303 13578 856
rect 13746 303 13762 856
rect 13930 303 13946 856
rect 14114 303 14130 856
rect 14298 303 14314 856
rect 14574 303 14590 856
rect 14758 303 14774 856
rect 14942 303 14958 856
rect 15126 303 15142 856
rect 15310 303 15326 856
rect 15494 303 15510 856
rect 15678 303 15694 856
rect 15862 303 15878 856
rect 16046 303 16062 856
rect 16230 303 16246 856
rect 16414 303 16430 856
rect 16598 303 16614 856
rect 16874 303 16890 856
rect 17058 303 17074 856
rect 17242 303 17258 856
rect 17426 303 17442 856
rect 17610 303 17626 856
rect 17794 303 17810 856
rect 17978 303 17994 856
rect 18162 303 18178 856
rect 18346 303 18362 856
rect 18530 303 18546 856
rect 18714 303 18730 856
rect 18898 303 18914 856
rect 19082 303 19098 856
rect 19358 303 19374 856
rect 19542 303 19558 856
rect 19726 303 19742 856
rect 19910 303 19926 856
rect 20094 303 20110 856
rect 20278 303 20294 856
rect 20462 303 20478 856
rect 20646 303 20662 856
rect 20830 303 20846 856
rect 21014 303 21030 856
rect 21198 303 21214 856
rect 21382 303 21398 856
rect 21658 303 21674 856
rect 21842 303 21858 856
rect 22026 303 22042 856
rect 22210 303 22226 856
rect 22394 303 22410 856
rect 22578 303 22594 856
rect 22762 303 22778 856
rect 22946 303 22962 856
rect 23130 303 23146 856
rect 23314 303 23330 856
rect 23498 303 23514 856
rect 23682 303 23698 856
rect 23866 303 23882 856
rect 24142 303 24158 856
rect 24326 303 24342 856
rect 24510 303 24526 856
rect 24694 303 24710 856
rect 24878 303 24894 856
rect 25062 303 25078 856
rect 25246 303 25262 856
rect 25430 303 25446 856
rect 25614 303 25630 856
rect 25798 303 25814 856
rect 25982 303 25998 856
rect 26166 303 26182 856
rect 26442 303 26458 856
rect 26626 303 26642 856
rect 26810 303 26826 856
rect 26994 303 27010 856
rect 27178 303 27194 856
rect 27362 303 27378 856
rect 27546 303 27562 856
rect 27730 303 27746 856
rect 27914 303 27930 856
rect 28098 303 28114 856
rect 28282 303 28298 856
rect 28466 303 28482 856
rect 28650 303 28666 856
rect 28926 303 28942 856
rect 29110 303 29126 856
rect 29294 303 29310 856
rect 29478 303 29494 856
rect 29662 303 29678 856
rect 29846 303 29862 856
rect 30030 303 30046 856
rect 30214 303 30230 856
rect 30398 303 30414 856
rect 30582 303 30598 856
rect 30766 303 30782 856
rect 30950 303 30966 856
rect 31226 303 31242 856
rect 31410 303 31426 856
rect 31594 303 31610 856
rect 31778 303 31794 856
rect 31962 303 31978 856
rect 32146 303 32162 856
rect 32330 303 32346 856
rect 32514 303 32530 856
rect 32698 303 32714 856
rect 32882 303 32898 856
rect 33066 303 33082 856
rect 33250 303 33266 856
rect 33434 303 33450 856
rect 33710 303 33726 856
rect 33894 303 33910 856
rect 34078 303 34094 856
rect 34262 303 34278 856
rect 34446 303 34462 856
rect 34630 303 34646 856
rect 34814 303 34830 856
rect 34998 303 35014 856
rect 35182 303 35198 856
rect 35366 303 35382 856
rect 35550 303 35566 856
rect 35734 303 35750 856
rect 36010 303 36026 856
rect 36194 303 36210 856
rect 36378 303 36394 856
rect 36562 303 36578 856
rect 36746 303 36762 856
rect 36930 303 36946 856
rect 37114 303 37130 856
rect 37298 303 37314 856
rect 37482 303 37498 856
rect 37666 303 37682 856
rect 37850 303 37866 856
rect 38034 303 38050 856
rect 38218 303 38234 856
rect 38494 303 38510 856
rect 38678 303 38694 856
rect 38862 303 38878 856
rect 39046 303 39062 856
rect 39230 303 39246 856
rect 39414 303 39430 856
rect 39598 303 39614 856
rect 39782 303 39798 856
rect 39966 303 39982 856
rect 40150 303 40166 856
rect 40334 303 40350 856
rect 40518 303 40534 856
rect 40794 303 40810 856
rect 40978 303 40994 856
rect 41162 303 41178 856
rect 41346 303 41362 856
rect 41530 303 41546 856
rect 41714 303 41730 856
rect 41898 303 41914 856
rect 42082 303 42098 856
rect 42266 303 42282 856
rect 42450 303 42466 856
rect 42634 303 42650 856
rect 42818 303 42834 856
rect 43002 303 43018 856
rect 43278 303 43294 856
rect 43462 303 43478 856
rect 43646 303 43662 856
rect 43830 303 43846 856
rect 44014 303 44030 856
rect 44198 303 44214 856
rect 44382 303 44398 856
rect 44566 303 44582 856
rect 44750 303 44766 856
rect 44934 303 44950 856
rect 45118 303 45134 856
rect 45302 303 45318 856
rect 45578 303 45594 856
rect 45762 303 45778 856
rect 45946 303 45962 856
rect 46130 303 46146 856
rect 46314 303 46330 856
rect 46498 303 46514 856
rect 46682 303 46698 856
rect 46866 303 46882 856
rect 47050 303 47066 856
rect 47234 303 47250 856
rect 47418 303 47434 856
rect 47602 303 47618 856
rect 47786 303 47802 856
rect 48062 303 48078 856
rect 48246 303 48262 856
rect 48430 303 48446 856
rect 48614 303 48630 856
rect 48798 303 48814 856
rect 48982 303 48998 856
rect 49166 303 49182 856
rect 49350 303 49366 856
rect 49534 303 49550 856
rect 49718 303 49734 856
rect 49902 303 49918 856
rect 50086 303 50102 856
rect 50362 303 50378 856
rect 50546 303 50562 856
rect 50730 303 50746 856
rect 50914 303 50930 856
rect 51098 303 51114 856
rect 51282 303 51298 856
rect 51466 303 51482 856
rect 51650 303 51666 856
rect 51834 303 51850 856
rect 52018 303 52034 856
rect 52202 303 52218 856
rect 52386 303 52402 856
rect 52570 303 52586 856
rect 52846 303 52862 856
rect 53030 303 53046 856
rect 53214 303 53230 856
rect 53398 303 53414 856
rect 53582 303 53598 856
rect 53766 303 53782 856
rect 53950 303 53966 856
rect 54134 303 54150 856
rect 54318 303 54334 856
rect 54502 303 54518 856
rect 54686 303 54702 856
rect 54870 303 54886 856
rect 55146 303 55162 856
rect 55330 303 55346 856
rect 55514 303 55530 856
rect 55698 303 55714 856
rect 55882 303 55898 856
rect 56066 303 56082 856
rect 56250 303 56266 856
rect 56434 303 56450 856
rect 56618 303 56634 856
rect 56802 303 56818 856
rect 56986 303 57002 856
rect 57170 303 57186 856
rect 57354 303 57370 856
rect 57630 303 57646 856
rect 57814 303 57830 856
rect 57998 303 58014 856
rect 58182 303 58198 856
rect 58366 303 58382 856
rect 58550 303 58566 856
rect 58734 303 58750 856
rect 58918 303 58934 856
rect 59102 303 59118 856
rect 59286 303 59302 856
rect 59470 303 59486 856
rect 59654 303 59670 856
rect 59838 303 59854 856
rect 60114 303 60130 856
rect 60298 303 60314 856
rect 60482 303 60498 856
rect 60666 303 60682 856
rect 60850 303 60866 856
rect 61034 303 61050 856
rect 61218 303 61234 856
rect 61402 303 61418 856
rect 61586 303 61602 856
rect 61770 303 61786 856
rect 61954 303 61970 856
rect 62138 303 62154 856
rect 62414 303 62430 856
rect 62598 303 62614 856
rect 62782 303 62798 856
rect 62966 303 62982 856
rect 63150 303 63166 856
rect 63334 303 63350 856
rect 63518 303 63534 856
rect 63702 303 63718 856
rect 63886 303 63902 856
rect 64070 303 64086 856
rect 64254 303 64270 856
rect 64438 303 64454 856
rect 64622 303 64638 856
rect 64898 303 64914 856
rect 65082 303 65098 856
rect 65266 303 65282 856
rect 65450 303 65466 856
rect 65634 303 65650 856
rect 65818 303 65834 856
rect 66002 303 66018 856
rect 66186 303 66202 856
rect 66370 303 66386 856
rect 66554 303 66570 856
rect 66738 303 66754 856
rect 66922 303 66938 856
rect 67198 303 67214 856
rect 67382 303 67398 856
rect 67566 303 67582 856
rect 67750 303 67766 856
rect 67934 303 67950 856
rect 68118 303 68134 856
rect 68302 303 68318 856
rect 68486 303 68502 856
rect 68670 303 68686 856
rect 68854 303 68870 856
rect 69038 303 69054 856
rect 69222 303 69238 856
rect 69406 303 69422 856
rect 69682 303 69698 856
rect 69866 303 69882 856
rect 70050 303 70066 856
rect 70234 303 70250 856
rect 70418 303 70434 856
rect 70602 303 70618 856
rect 70786 303 70802 856
rect 70970 303 70986 856
rect 71154 303 71170 856
rect 71338 303 71354 856
rect 71522 303 71538 856
rect 71706 303 71722 856
rect 71982 303 71998 856
rect 72166 303 72182 856
rect 72350 303 72366 856
rect 72534 303 72550 856
rect 72718 303 72734 856
rect 72902 303 72918 856
rect 73086 303 73102 856
rect 73270 303 73286 856
rect 73454 303 73470 856
rect 73638 303 73654 856
rect 73822 303 73838 856
rect 74006 303 74022 856
rect 74190 303 74206 856
rect 74466 303 74482 856
rect 74650 303 74666 856
rect 74834 303 74850 856
rect 75018 303 75034 856
rect 75202 303 75218 856
rect 75386 303 75402 856
rect 75570 303 75586 856
rect 75754 303 75770 856
rect 75938 303 75954 856
rect 76122 303 76138 856
rect 76306 303 76322 856
rect 76490 303 76506 856
rect 76766 303 76782 856
rect 76950 303 76966 856
rect 77134 303 77150 856
rect 77318 303 77334 856
rect 77502 303 77518 856
rect 77686 303 77702 856
rect 77870 303 77886 856
rect 78054 303 78070 856
rect 78238 303 78254 856
rect 78422 303 78438 856
rect 78606 303 78622 856
rect 78790 303 78806 856
rect 78974 303 78990 856
rect 79250 303 79266 856
rect 79434 303 79450 856
rect 79618 303 79634 856
rect 79802 303 79818 856
rect 79986 303 80002 856
rect 80170 303 80186 856
rect 80354 303 80370 856
rect 80538 303 80554 856
rect 80722 303 80738 856
rect 80906 303 80922 856
rect 81090 303 81106 856
rect 81274 303 81290 856
rect 81550 303 81566 856
rect 81734 303 81750 856
rect 81918 303 81934 856
rect 82102 303 82118 856
rect 82286 303 82302 856
rect 82470 303 82486 856
rect 82654 303 82670 856
rect 82838 303 82854 856
rect 83022 303 83038 856
rect 83206 303 83222 856
rect 83390 303 83406 856
rect 83574 303 83590 856
rect 83758 303 83774 856
rect 84034 303 84050 856
rect 84218 303 84234 856
rect 84402 303 84418 856
rect 84586 303 84602 856
rect 84770 303 84786 856
rect 84954 303 84970 856
rect 85138 303 85154 856
rect 85322 303 85338 856
rect 85506 303 85522 856
rect 85690 303 85706 856
rect 85874 303 85890 856
rect 86058 303 86074 856
rect 86334 303 86350 856
rect 86518 303 86534 856
rect 86702 303 86718 856
rect 86886 303 86902 856
rect 87070 303 87086 856
rect 87254 303 87270 856
rect 87438 303 87454 856
rect 87622 303 87638 856
rect 87806 303 87822 856
rect 87990 303 88006 856
rect 88174 303 88190 856
rect 88358 303 88374 856
rect 88542 303 88558 856
rect 88818 303 88834 856
rect 89002 303 89018 856
rect 89186 303 89202 856
rect 89370 303 89386 856
rect 89554 303 89570 856
rect 89738 303 89754 856
rect 89922 303 89938 856
rect 90106 303 90122 856
rect 90290 303 90306 856
rect 90474 303 90490 856
rect 90658 303 90674 856
rect 90842 303 90858 856
rect 91118 303 91134 856
rect 91302 303 91318 856
rect 91486 303 91502 856
rect 91670 303 91686 856
rect 91854 303 91870 856
rect 92038 303 92054 856
rect 92222 303 92238 856
rect 92406 303 92422 856
rect 92590 303 92606 856
rect 92774 303 92790 856
rect 92958 303 92974 856
rect 93142 303 93158 856
rect 93326 303 93342 856
rect 93602 303 93618 856
rect 93786 303 93802 856
rect 93970 303 93986 856
rect 94154 303 94170 856
rect 94338 303 94354 856
rect 94522 303 94538 856
rect 94706 303 94722 856
rect 94890 303 94906 856
rect 95074 303 95090 856
rect 95258 303 95274 856
rect 95442 303 95458 856
rect 95626 303 95642 856
rect 95902 303 95918 856
rect 96086 303 96102 856
rect 96270 303 96286 856
rect 96454 303 96470 856
rect 96638 303 96654 856
rect 96822 303 96838 856
rect 97006 303 97022 856
rect 97190 303 97206 856
rect 97374 303 97390 856
rect 97558 303 97574 856
rect 97742 303 97758 856
rect 97926 303 97942 856
rect 98110 303 98126 856
rect 98386 303 98402 856
rect 98570 303 98586 856
rect 98754 303 98770 856
rect 98938 303 98954 856
rect 99122 303 99138 856
rect 99306 303 99322 856
rect 99490 303 99506 856
rect 99674 303 99690 856
rect 99858 303 99874 856
rect 100042 303 100058 856
rect 100226 303 100242 856
rect 100410 303 100426 856
rect 100686 303 100702 856
rect 100870 303 100886 856
rect 101054 303 101070 856
rect 101238 303 101254 856
rect 101422 303 101438 856
rect 101606 303 101622 856
rect 101790 303 101806 856
rect 101974 303 101990 856
rect 102158 303 102174 856
rect 102342 303 102358 856
rect 102526 303 102542 856
rect 102710 303 102726 856
rect 102894 303 102910 856
rect 103170 303 103186 856
rect 103354 303 103370 856
rect 103538 303 103554 856
rect 103722 303 103738 856
rect 103906 303 103922 856
rect 104090 303 104106 856
rect 104274 303 104290 856
rect 104458 303 104474 856
rect 104642 303 104658 856
rect 104826 303 104842 856
rect 105010 303 105026 856
rect 105194 303 105210 856
rect 105470 303 105486 856
rect 105654 303 105670 856
rect 105838 303 105854 856
rect 106022 303 106038 856
rect 106206 303 106222 856
rect 106390 303 106406 856
rect 106574 303 106590 856
rect 106758 303 106774 856
rect 106942 303 106958 856
rect 107126 303 107142 856
rect 107310 303 107326 856
rect 107494 303 107510 856
rect 107678 303 107694 856
rect 107954 303 107970 856
rect 108138 303 108154 856
rect 108322 303 108338 856
rect 108506 303 108522 856
rect 108690 303 108706 856
rect 108874 303 108890 856
rect 109058 303 109074 856
rect 109242 303 109258 856
rect 109426 303 109442 856
rect 109610 303 109626 856
rect 109794 303 109810 856
rect 109978 303 109994 856
rect 110254 303 110270 856
rect 110438 303 110454 856
rect 110622 303 110638 856
rect 110806 303 110822 856
rect 110990 303 111006 856
rect 111174 303 111190 856
rect 111358 303 111374 856
rect 111542 303 111558 856
rect 111726 303 111742 856
rect 111910 303 111926 856
rect 112094 303 112110 856
rect 112278 303 112294 856
rect 112462 303 112478 856
rect 112738 303 112754 856
rect 112922 303 112938 856
rect 113106 303 113122 856
rect 113290 303 113306 856
rect 113474 303 113490 856
rect 113658 303 113674 856
rect 113842 303 113858 856
rect 114026 303 114042 856
rect 114210 303 114226 856
rect 114394 303 114410 856
rect 114578 303 114594 856
rect 114762 303 114778 856
rect 115038 303 115054 856
rect 115222 303 115238 856
rect 115406 303 115422 856
rect 115590 303 115606 856
rect 115774 303 115790 856
rect 115958 303 115974 856
rect 116142 303 116158 856
rect 116326 303 116342 856
rect 116510 303 116526 856
rect 116694 303 116710 856
rect 116878 303 116894 856
rect 117062 303 117078 856
rect 117246 303 117262 856
rect 117522 303 117538 856
rect 117706 303 117722 856
rect 117890 303 117906 856
rect 118074 303 118090 856
rect 118258 303 118274 856
rect 118442 303 118458 856
rect 118626 303 118642 856
rect 118810 303 118826 856
rect 118994 303 119010 856
rect 119178 303 119194 856
rect 119362 303 119378 856
rect 119546 303 119562 856
<< obsm3 >>
rect 13 307 119311 119713
<< metal4 >>
rect 4208 2128 4528 119728
rect 19568 2128 19888 119728
rect 34928 2128 35248 119728
rect 50288 2128 50608 119728
rect 65648 2128 65968 119728
rect 81008 2128 81328 119728
rect 96368 2128 96688 119728
rect 111728 2128 112048 119728
<< obsm4 >>
rect 1899 2048 4128 119101
rect 4608 2048 19488 119101
rect 19968 2048 34848 119101
rect 35328 2048 50208 119101
rect 50688 2048 65568 119101
rect 66048 2048 80928 119101
rect 81408 2048 96288 119101
rect 96768 2048 111648 119101
rect 112128 2048 117517 119101
rect 1899 307 117517 2048
<< labels >>
rlabel metal2 s 71410 121102 71466 121902 6 dram_addr0[0]
port 1 nsew signal output
rlabel metal2 s 73802 121102 73858 121902 6 dram_addr0[1]
port 2 nsew signal output
rlabel metal2 s 76286 121102 76342 121902 6 dram_addr0[2]
port 3 nsew signal output
rlabel metal2 s 78678 121102 78734 121902 6 dram_addr0[3]
port 4 nsew signal output
rlabel metal2 s 81162 121102 81218 121902 6 dram_addr0[4]
port 5 nsew signal output
rlabel metal2 s 82910 121102 82966 121902 6 dram_addr0[5]
port 6 nsew signal output
rlabel metal2 s 84750 121102 84806 121902 6 dram_addr0[6]
port 7 nsew signal output
rlabel metal2 s 86590 121102 86646 121902 6 dram_addr0[7]
port 8 nsew signal output
rlabel metal2 s 88430 121102 88486 121902 6 dram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 69570 121102 69626 121902 6 dram_clk0
port 10 nsew signal output
rlabel metal2 s 70214 121102 70270 121902 6 dram_csb0
port 11 nsew signal output
rlabel metal2 s 71962 121102 72018 121902 6 dram_din0[0]
port 12 nsew signal output
rlabel metal2 s 91466 121102 91522 121902 6 dram_din0[10]
port 13 nsew signal output
rlabel metal2 s 92662 121102 92718 121902 6 dram_din0[11]
port 14 nsew signal output
rlabel metal2 s 93858 121102 93914 121902 6 dram_din0[12]
port 15 nsew signal output
rlabel metal2 s 95146 121102 95202 121902 6 dram_din0[13]
port 16 nsew signal output
rlabel metal2 s 96342 121102 96398 121902 6 dram_din0[14]
port 17 nsew signal output
rlabel metal2 s 97538 121102 97594 121902 6 dram_din0[15]
port 18 nsew signal output
rlabel metal2 s 98734 121102 98790 121902 6 dram_din0[16]
port 19 nsew signal output
rlabel metal2 s 99930 121102 99986 121902 6 dram_din0[17]
port 20 nsew signal output
rlabel metal2 s 101218 121102 101274 121902 6 dram_din0[18]
port 21 nsew signal output
rlabel metal2 s 102414 121102 102470 121902 6 dram_din0[19]
port 22 nsew signal output
rlabel metal2 s 74446 121102 74502 121902 6 dram_din0[1]
port 23 nsew signal output
rlabel metal2 s 103610 121102 103666 121902 6 dram_din0[20]
port 24 nsew signal output
rlabel metal2 s 104806 121102 104862 121902 6 dram_din0[21]
port 25 nsew signal output
rlabel metal2 s 106002 121102 106058 121902 6 dram_din0[22]
port 26 nsew signal output
rlabel metal2 s 107290 121102 107346 121902 6 dram_din0[23]
port 27 nsew signal output
rlabel metal2 s 108486 121102 108542 121902 6 dram_din0[24]
port 28 nsew signal output
rlabel metal2 s 109682 121102 109738 121902 6 dram_din0[25]
port 29 nsew signal output
rlabel metal2 s 110878 121102 110934 121902 6 dram_din0[26]
port 30 nsew signal output
rlabel metal2 s 112166 121102 112222 121902 6 dram_din0[27]
port 31 nsew signal output
rlabel metal2 s 113362 121102 113418 121902 6 dram_din0[28]
port 32 nsew signal output
rlabel metal2 s 114558 121102 114614 121902 6 dram_din0[29]
port 33 nsew signal output
rlabel metal2 s 76838 121102 76894 121902 6 dram_din0[2]
port 34 nsew signal output
rlabel metal2 s 115754 121102 115810 121902 6 dram_din0[30]
port 35 nsew signal output
rlabel metal2 s 116950 121102 117006 121902 6 dram_din0[31]
port 36 nsew signal output
rlabel metal2 s 79322 121102 79378 121902 6 dram_din0[3]
port 37 nsew signal output
rlabel metal2 s 81714 121102 81770 121902 6 dram_din0[4]
port 38 nsew signal output
rlabel metal2 s 83554 121102 83610 121902 6 dram_din0[5]
port 39 nsew signal output
rlabel metal2 s 85394 121102 85450 121902 6 dram_din0[6]
port 40 nsew signal output
rlabel metal2 s 87234 121102 87290 121902 6 dram_din0[7]
port 41 nsew signal output
rlabel metal2 s 88982 121102 89038 121902 6 dram_din0[8]
port 42 nsew signal output
rlabel metal2 s 90270 121102 90326 121902 6 dram_din0[9]
port 43 nsew signal output
rlabel metal2 s 72606 121102 72662 121902 6 dram_dout0[0]
port 44 nsew signal input
rlabel metal2 s 92018 121102 92074 121902 6 dram_dout0[10]
port 45 nsew signal input
rlabel metal2 s 93306 121102 93362 121902 6 dram_dout0[11]
port 46 nsew signal input
rlabel metal2 s 94502 121102 94558 121902 6 dram_dout0[12]
port 47 nsew signal input
rlabel metal2 s 95698 121102 95754 121902 6 dram_dout0[13]
port 48 nsew signal input
rlabel metal2 s 96894 121102 96950 121902 6 dram_dout0[14]
port 49 nsew signal input
rlabel metal2 s 98182 121102 98238 121902 6 dram_dout0[15]
port 50 nsew signal input
rlabel metal2 s 99378 121102 99434 121902 6 dram_dout0[16]
port 51 nsew signal input
rlabel metal2 s 100574 121102 100630 121902 6 dram_dout0[17]
port 52 nsew signal input
rlabel metal2 s 101770 121102 101826 121902 6 dram_dout0[18]
port 53 nsew signal input
rlabel metal2 s 102966 121102 103022 121902 6 dram_dout0[19]
port 54 nsew signal input
rlabel metal2 s 74998 121102 75054 121902 6 dram_dout0[1]
port 55 nsew signal input
rlabel metal2 s 104254 121102 104310 121902 6 dram_dout0[20]
port 56 nsew signal input
rlabel metal2 s 105450 121102 105506 121902 6 dram_dout0[21]
port 57 nsew signal input
rlabel metal2 s 106646 121102 106702 121902 6 dram_dout0[22]
port 58 nsew signal input
rlabel metal2 s 107842 121102 107898 121902 6 dram_dout0[23]
port 59 nsew signal input
rlabel metal2 s 109130 121102 109186 121902 6 dram_dout0[24]
port 60 nsew signal input
rlabel metal2 s 110326 121102 110382 121902 6 dram_dout0[25]
port 61 nsew signal input
rlabel metal2 s 111522 121102 111578 121902 6 dram_dout0[26]
port 62 nsew signal input
rlabel metal2 s 112718 121102 112774 121902 6 dram_dout0[27]
port 63 nsew signal input
rlabel metal2 s 113914 121102 113970 121902 6 dram_dout0[28]
port 64 nsew signal input
rlabel metal2 s 115202 121102 115258 121902 6 dram_dout0[29]
port 65 nsew signal input
rlabel metal2 s 77482 121102 77538 121902 6 dram_dout0[2]
port 66 nsew signal input
rlabel metal2 s 116398 121102 116454 121902 6 dram_dout0[30]
port 67 nsew signal input
rlabel metal2 s 117594 121102 117650 121902 6 dram_dout0[31]
port 68 nsew signal input
rlabel metal2 s 79874 121102 79930 121902 6 dram_dout0[3]
port 69 nsew signal input
rlabel metal2 s 82358 121102 82414 121902 6 dram_dout0[4]
port 70 nsew signal input
rlabel metal2 s 84198 121102 84254 121902 6 dram_dout0[5]
port 71 nsew signal input
rlabel metal2 s 85946 121102 86002 121902 6 dram_dout0[6]
port 72 nsew signal input
rlabel metal2 s 87786 121102 87842 121902 6 dram_dout0[7]
port 73 nsew signal input
rlabel metal2 s 89626 121102 89682 121902 6 dram_dout0[8]
port 74 nsew signal input
rlabel metal2 s 90822 121102 90878 121902 6 dram_dout0[9]
port 75 nsew signal input
rlabel metal2 s 70766 121102 70822 121902 6 dram_web0
port 76 nsew signal output
rlabel metal2 s 73250 121102 73306 121902 6 dram_wmask0[0]
port 77 nsew signal output
rlabel metal2 s 75642 121102 75698 121902 6 dram_wmask0[1]
port 78 nsew signal output
rlabel metal2 s 78034 121102 78090 121902 6 dram_wmask0[2]
port 79 nsew signal output
rlabel metal2 s 80518 121102 80574 121902 6 dram_wmask0[3]
port 80 nsew signal output
rlabel metal2 s 294 121102 350 121902 6 io_in[0]
port 81 nsew signal input
rlabel metal2 s 18510 121102 18566 121902 6 io_in[10]
port 82 nsew signal input
rlabel metal2 s 20350 121102 20406 121902 6 io_in[11]
port 83 nsew signal input
rlabel metal2 s 22098 121102 22154 121902 6 io_in[12]
port 84 nsew signal input
rlabel metal2 s 23938 121102 23994 121902 6 io_in[13]
port 85 nsew signal input
rlabel metal2 s 25778 121102 25834 121902 6 io_in[14]
port 86 nsew signal input
rlabel metal2 s 27618 121102 27674 121902 6 io_in[15]
port 87 nsew signal input
rlabel metal2 s 29458 121102 29514 121902 6 io_in[16]
port 88 nsew signal input
rlabel metal2 s 31298 121102 31354 121902 6 io_in[17]
port 89 nsew signal input
rlabel metal2 s 33046 121102 33102 121902 6 io_in[18]
port 90 nsew signal input
rlabel metal2 s 34886 121102 34942 121902 6 io_in[19]
port 91 nsew signal input
rlabel metal2 s 2042 121102 2098 121902 6 io_in[1]
port 92 nsew signal input
rlabel metal2 s 36726 121102 36782 121902 6 io_in[20]
port 93 nsew signal input
rlabel metal2 s 38566 121102 38622 121902 6 io_in[21]
port 94 nsew signal input
rlabel metal2 s 40406 121102 40462 121902 6 io_in[22]
port 95 nsew signal input
rlabel metal2 s 42246 121102 42302 121902 6 io_in[23]
port 96 nsew signal input
rlabel metal2 s 43994 121102 44050 121902 6 io_in[24]
port 97 nsew signal input
rlabel metal2 s 45834 121102 45890 121902 6 io_in[25]
port 98 nsew signal input
rlabel metal2 s 47674 121102 47730 121902 6 io_in[26]
port 99 nsew signal input
rlabel metal2 s 49514 121102 49570 121902 6 io_in[27]
port 100 nsew signal input
rlabel metal2 s 51354 121102 51410 121902 6 io_in[28]
port 101 nsew signal input
rlabel metal2 s 53102 121102 53158 121902 6 io_in[29]
port 102 nsew signal input
rlabel metal2 s 3882 121102 3938 121902 6 io_in[2]
port 103 nsew signal input
rlabel metal2 s 54942 121102 54998 121902 6 io_in[30]
port 104 nsew signal input
rlabel metal2 s 56782 121102 56838 121902 6 io_in[31]
port 105 nsew signal input
rlabel metal2 s 58622 121102 58678 121902 6 io_in[32]
port 106 nsew signal input
rlabel metal2 s 60462 121102 60518 121902 6 io_in[33]
port 107 nsew signal input
rlabel metal2 s 62302 121102 62358 121902 6 io_in[34]
port 108 nsew signal input
rlabel metal2 s 64050 121102 64106 121902 6 io_in[35]
port 109 nsew signal input
rlabel metal2 s 65890 121102 65946 121902 6 io_in[36]
port 110 nsew signal input
rlabel metal2 s 67730 121102 67786 121902 6 io_in[37]
port 111 nsew signal input
rlabel metal2 s 5722 121102 5778 121902 6 io_in[3]
port 112 nsew signal input
rlabel metal2 s 7562 121102 7618 121902 6 io_in[4]
port 113 nsew signal input
rlabel metal2 s 9402 121102 9458 121902 6 io_in[5]
port 114 nsew signal input
rlabel metal2 s 11150 121102 11206 121902 6 io_in[6]
port 115 nsew signal input
rlabel metal2 s 12990 121102 13046 121902 6 io_in[7]
port 116 nsew signal input
rlabel metal2 s 14830 121102 14886 121902 6 io_in[8]
port 117 nsew signal input
rlabel metal2 s 16670 121102 16726 121902 6 io_in[9]
port 118 nsew signal input
rlabel metal2 s 846 121102 902 121902 6 io_oeb[0]
port 119 nsew signal output
rlabel metal2 s 19062 121102 19118 121902 6 io_oeb[10]
port 120 nsew signal output
rlabel metal2 s 20902 121102 20958 121902 6 io_oeb[11]
port 121 nsew signal output
rlabel metal2 s 22742 121102 22798 121902 6 io_oeb[12]
port 122 nsew signal output
rlabel metal2 s 24582 121102 24638 121902 6 io_oeb[13]
port 123 nsew signal output
rlabel metal2 s 26422 121102 26478 121902 6 io_oeb[14]
port 124 nsew signal output
rlabel metal2 s 28262 121102 28318 121902 6 io_oeb[15]
port 125 nsew signal output
rlabel metal2 s 30010 121102 30066 121902 6 io_oeb[16]
port 126 nsew signal output
rlabel metal2 s 31850 121102 31906 121902 6 io_oeb[17]
port 127 nsew signal output
rlabel metal2 s 33690 121102 33746 121902 6 io_oeb[18]
port 128 nsew signal output
rlabel metal2 s 35530 121102 35586 121902 6 io_oeb[19]
port 129 nsew signal output
rlabel metal2 s 2686 121102 2742 121902 6 io_oeb[1]
port 130 nsew signal output
rlabel metal2 s 37370 121102 37426 121902 6 io_oeb[20]
port 131 nsew signal output
rlabel metal2 s 39118 121102 39174 121902 6 io_oeb[21]
port 132 nsew signal output
rlabel metal2 s 40958 121102 41014 121902 6 io_oeb[22]
port 133 nsew signal output
rlabel metal2 s 42798 121102 42854 121902 6 io_oeb[23]
port 134 nsew signal output
rlabel metal2 s 44638 121102 44694 121902 6 io_oeb[24]
port 135 nsew signal output
rlabel metal2 s 46478 121102 46534 121902 6 io_oeb[25]
port 136 nsew signal output
rlabel metal2 s 48318 121102 48374 121902 6 io_oeb[26]
port 137 nsew signal output
rlabel metal2 s 50066 121102 50122 121902 6 io_oeb[27]
port 138 nsew signal output
rlabel metal2 s 51906 121102 51962 121902 6 io_oeb[28]
port 139 nsew signal output
rlabel metal2 s 53746 121102 53802 121902 6 io_oeb[29]
port 140 nsew signal output
rlabel metal2 s 4526 121102 4582 121902 6 io_oeb[2]
port 141 nsew signal output
rlabel metal2 s 55586 121102 55642 121902 6 io_oeb[30]
port 142 nsew signal output
rlabel metal2 s 57426 121102 57482 121902 6 io_oeb[31]
port 143 nsew signal output
rlabel metal2 s 59266 121102 59322 121902 6 io_oeb[32]
port 144 nsew signal output
rlabel metal2 s 61014 121102 61070 121902 6 io_oeb[33]
port 145 nsew signal output
rlabel metal2 s 62854 121102 62910 121902 6 io_oeb[34]
port 146 nsew signal output
rlabel metal2 s 64694 121102 64750 121902 6 io_oeb[35]
port 147 nsew signal output
rlabel metal2 s 66534 121102 66590 121902 6 io_oeb[36]
port 148 nsew signal output
rlabel metal2 s 68374 121102 68430 121902 6 io_oeb[37]
port 149 nsew signal output
rlabel metal2 s 6366 121102 6422 121902 6 io_oeb[3]
port 150 nsew signal output
rlabel metal2 s 8114 121102 8170 121902 6 io_oeb[4]
port 151 nsew signal output
rlabel metal2 s 9954 121102 10010 121902 6 io_oeb[5]
port 152 nsew signal output
rlabel metal2 s 11794 121102 11850 121902 6 io_oeb[6]
port 153 nsew signal output
rlabel metal2 s 13634 121102 13690 121902 6 io_oeb[7]
port 154 nsew signal output
rlabel metal2 s 15474 121102 15530 121902 6 io_oeb[8]
port 155 nsew signal output
rlabel metal2 s 17314 121102 17370 121902 6 io_oeb[9]
port 156 nsew signal output
rlabel metal2 s 1490 121102 1546 121902 6 io_out[0]
port 157 nsew signal output
rlabel metal2 s 19706 121102 19762 121902 6 io_out[10]
port 158 nsew signal output
rlabel metal2 s 21546 121102 21602 121902 6 io_out[11]
port 159 nsew signal output
rlabel metal2 s 23386 121102 23442 121902 6 io_out[12]
port 160 nsew signal output
rlabel metal2 s 25134 121102 25190 121902 6 io_out[13]
port 161 nsew signal output
rlabel metal2 s 26974 121102 27030 121902 6 io_out[14]
port 162 nsew signal output
rlabel metal2 s 28814 121102 28870 121902 6 io_out[15]
port 163 nsew signal output
rlabel metal2 s 30654 121102 30710 121902 6 io_out[16]
port 164 nsew signal output
rlabel metal2 s 32494 121102 32550 121902 6 io_out[17]
port 165 nsew signal output
rlabel metal2 s 34334 121102 34390 121902 6 io_out[18]
port 166 nsew signal output
rlabel metal2 s 36082 121102 36138 121902 6 io_out[19]
port 167 nsew signal output
rlabel metal2 s 3330 121102 3386 121902 6 io_out[1]
port 168 nsew signal output
rlabel metal2 s 37922 121102 37978 121902 6 io_out[20]
port 169 nsew signal output
rlabel metal2 s 39762 121102 39818 121902 6 io_out[21]
port 170 nsew signal output
rlabel metal2 s 41602 121102 41658 121902 6 io_out[22]
port 171 nsew signal output
rlabel metal2 s 43442 121102 43498 121902 6 io_out[23]
port 172 nsew signal output
rlabel metal2 s 45282 121102 45338 121902 6 io_out[24]
port 173 nsew signal output
rlabel metal2 s 47030 121102 47086 121902 6 io_out[25]
port 174 nsew signal output
rlabel metal2 s 48870 121102 48926 121902 6 io_out[26]
port 175 nsew signal output
rlabel metal2 s 50710 121102 50766 121902 6 io_out[27]
port 176 nsew signal output
rlabel metal2 s 52550 121102 52606 121902 6 io_out[28]
port 177 nsew signal output
rlabel metal2 s 54390 121102 54446 121902 6 io_out[29]
port 178 nsew signal output
rlabel metal2 s 5078 121102 5134 121902 6 io_out[2]
port 179 nsew signal output
rlabel metal2 s 56230 121102 56286 121902 6 io_out[30]
port 180 nsew signal output
rlabel metal2 s 57978 121102 58034 121902 6 io_out[31]
port 181 nsew signal output
rlabel metal2 s 59818 121102 59874 121902 6 io_out[32]
port 182 nsew signal output
rlabel metal2 s 61658 121102 61714 121902 6 io_out[33]
port 183 nsew signal output
rlabel metal2 s 63498 121102 63554 121902 6 io_out[34]
port 184 nsew signal output
rlabel metal2 s 65338 121102 65394 121902 6 io_out[35]
port 185 nsew signal output
rlabel metal2 s 67178 121102 67234 121902 6 io_out[36]
port 186 nsew signal output
rlabel metal2 s 68926 121102 68982 121902 6 io_out[37]
port 187 nsew signal output
rlabel metal2 s 6918 121102 6974 121902 6 io_out[3]
port 188 nsew signal output
rlabel metal2 s 8758 121102 8814 121902 6 io_out[4]
port 189 nsew signal output
rlabel metal2 s 10598 121102 10654 121902 6 io_out[5]
port 190 nsew signal output
rlabel metal2 s 12438 121102 12494 121902 6 io_out[6]
port 191 nsew signal output
rlabel metal2 s 14278 121102 14334 121902 6 io_out[7]
port 192 nsew signal output
rlabel metal2 s 16026 121102 16082 121902 6 io_out[8]
port 193 nsew signal output
rlabel metal2 s 17866 121102 17922 121902 6 io_out[9]
port 194 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 iram_addr0[0]
port 195 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 iram_addr0[1]
port 196 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 iram_addr0[2]
port 197 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 iram_addr0[3]
port 198 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 iram_addr0[4]
port 199 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 iram_addr0[5]
port 200 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 iram_addr0[6]
port 201 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 iram_addr0[7]
port 202 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 iram_addr0[8]
port 203 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 iram_clk0
port 204 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 iram_csb0
port 205 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 iram_din0[0]
port 206 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 iram_din0[10]
port 207 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 iram_din0[11]
port 208 nsew signal output
rlabel metal2 s 112626 0 112682 800 6 iram_din0[12]
port 209 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 iram_din0[13]
port 210 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 iram_din0[14]
port 211 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 iram_din0[15]
port 212 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 iram_din0[16]
port 213 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 iram_din0[17]
port 214 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 iram_din0[18]
port 215 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 iram_din0[19]
port 216 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 iram_din0[1]
port 217 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 iram_din0[20]
port 218 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 iram_din0[21]
port 219 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 iram_din0[22]
port 220 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 iram_din0[23]
port 221 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 iram_din0[24]
port 222 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 iram_din0[25]
port 223 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 iram_din0[26]
port 224 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 iram_din0[27]
port 225 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 iram_din0[28]
port 226 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 iram_din0[29]
port 227 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 iram_din0[2]
port 228 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 iram_din0[30]
port 229 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 iram_din0[31]
port 230 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 iram_din0[3]
port 231 nsew signal output
rlabel metal2 s 109130 0 109186 800 6 iram_din0[4]
port 232 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 iram_din0[5]
port 233 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 iram_din0[6]
port 234 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 iram_din0[7]
port 235 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 iram_din0[8]
port 236 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 iram_din0[9]
port 237 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 iram_dout0[0]
port 238 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 iram_dout0[10]
port 239 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 iram_dout0[11]
port 240 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 iram_dout0[12]
port 241 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 iram_dout0[13]
port 242 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 iram_dout0[14]
port 243 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 iram_dout0[15]
port 244 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 iram_dout0[16]
port 245 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 iram_dout0[17]
port 246 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 iram_dout0[18]
port 247 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 iram_dout0[19]
port 248 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 iram_dout0[1]
port 249 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 iram_dout0[20]
port 250 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 iram_dout0[21]
port 251 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 iram_dout0[22]
port 252 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 iram_dout0[23]
port 253 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 iram_dout0[24]
port 254 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 iram_dout0[25]
port 255 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 iram_dout0[26]
port 256 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 iram_dout0[27]
port 257 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 iram_dout0[28]
port 258 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 iram_dout0[29]
port 259 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 iram_dout0[2]
port 260 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 iram_dout0[30]
port 261 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 iram_dout0[31]
port 262 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 iram_dout0[3]
port 263 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 iram_dout0[4]
port 264 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 iram_dout0[5]
port 265 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 iram_dout0[6]
port 266 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 iram_dout0[7]
port 267 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 iram_dout0[8]
port 268 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 iram_dout0[9]
port 269 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 iram_web0
port 270 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 iram_wmask0[0]
port 271 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 iram_wmask0[1]
port 272 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 iram_wmask0[2]
port 273 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 iram_wmask0[3]
port 274 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_in[0]
port 275 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[100]
port 276 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[101]
port 277 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[102]
port 278 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[103]
port 279 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[104]
port 280 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[105]
port 281 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[106]
port 282 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[107]
port 283 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[108]
port 284 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[109]
port 285 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[10]
port 286 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[110]
port 287 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[111]
port 288 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[112]
port 289 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[113]
port 290 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[114]
port 291 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[115]
port 292 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[116]
port 293 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_data_in[117]
port 294 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[118]
port 295 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[119]
port 296 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[11]
port 297 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_data_in[120]
port 298 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[121]
port 299 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_data_in[122]
port 300 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[123]
port 301 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[124]
port 302 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[125]
port 303 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[126]
port 304 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_data_in[127]
port 305 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[12]
port 306 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[13]
port 307 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[14]
port 308 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_data_in[15]
port 309 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[16]
port 310 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[17]
port 311 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[18]
port 312 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[19]
port 313 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[1]
port 314 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[20]
port 315 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[21]
port 316 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[22]
port 317 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[23]
port 318 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[24]
port 319 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[25]
port 320 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_data_in[26]
port 321 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[27]
port 322 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[28]
port 323 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[29]
port 324 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[2]
port 325 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[30]
port 326 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[31]
port 327 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[32]
port 328 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[33]
port 329 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[34]
port 330 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[35]
port 331 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[36]
port 332 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[37]
port 333 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[38]
port 334 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[39]
port 335 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[3]
port 336 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[40]
port 337 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[41]
port 338 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[42]
port 339 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_data_in[43]
port 340 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[44]
port 341 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[45]
port 342 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[46]
port 343 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[47]
port 344 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[48]
port 345 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[49]
port 346 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[4]
port 347 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[50]
port 348 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[51]
port 349 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[52]
port 350 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[53]
port 351 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[54]
port 352 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[55]
port 353 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[56]
port 354 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[57]
port 355 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[58]
port 356 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[59]
port 357 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[5]
port 358 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[60]
port 359 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[61]
port 360 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[62]
port 361 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[63]
port 362 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[64]
port 363 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[65]
port 364 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[66]
port 365 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[67]
port 366 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[68]
port 367 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[69]
port 368 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[6]
port 369 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_data_in[70]
port 370 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[71]
port 371 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[72]
port 372 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[73]
port 373 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_data_in[74]
port 374 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[75]
port 375 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[76]
port 376 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[77]
port 377 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[78]
port 378 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[79]
port 379 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[7]
port 380 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[80]
port 381 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[81]
port 382 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[82]
port 383 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[83]
port 384 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[84]
port 385 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[85]
port 386 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[86]
port 387 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[87]
port 388 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[88]
port 389 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[89]
port 390 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[8]
port 391 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[90]
port 392 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_data_in[91]
port 393 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[92]
port 394 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[93]
port 395 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[94]
port 396 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[95]
port 397 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[96]
port 398 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[97]
port 399 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_data_in[98]
port 400 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[99]
port 401 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[9]
port 402 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_data_out[0]
port 403 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[100]
port 404 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[101]
port 405 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[102]
port 406 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[103]
port 407 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[104]
port 408 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[105]
port 409 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[106]
port 410 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[107]
port 411 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[108]
port 412 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[109]
port 413 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[10]
port 414 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[110]
port 415 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[111]
port 416 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[112]
port 417 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[113]
port 418 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[114]
port 419 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[115]
port 420 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[116]
port 421 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[117]
port 422 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[118]
port 423 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[119]
port 424 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[11]
port 425 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 la_data_out[120]
port 426 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[121]
port 427 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[122]
port 428 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[123]
port 429 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[124]
port 430 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[125]
port 431 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[126]
port 432 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[127]
port 433 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[12]
port 434 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[13]
port 435 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[14]
port 436 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 la_data_out[15]
port 437 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[16]
port 438 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 la_data_out[17]
port 439 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[18]
port 440 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[19]
port 441 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[1]
port 442 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[20]
port 443 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[21]
port 444 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[22]
port 445 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[23]
port 446 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[24]
port 447 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[25]
port 448 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_data_out[26]
port 449 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[27]
port 450 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[28]
port 451 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[29]
port 452 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[2]
port 453 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[30]
port 454 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[31]
port 455 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[32]
port 456 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[33]
port 457 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[34]
port 458 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[35]
port 459 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[36]
port 460 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[37]
port 461 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[38]
port 462 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[39]
port 463 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[3]
port 464 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[40]
port 465 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[41]
port 466 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[42]
port 467 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_data_out[43]
port 468 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[44]
port 469 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 la_data_out[45]
port 470 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[46]
port 471 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 la_data_out[47]
port 472 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 la_data_out[48]
port 473 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[49]
port 474 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 la_data_out[4]
port 475 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[50]
port 476 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[51]
port 477 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[52]
port 478 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[53]
port 479 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[54]
port 480 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[55]
port 481 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[56]
port 482 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[57]
port 483 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 la_data_out[58]
port 484 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[59]
port 485 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[5]
port 486 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[60]
port 487 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[61]
port 488 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[62]
port 489 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[63]
port 490 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[64]
port 491 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[65]
port 492 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[66]
port 493 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[67]
port 494 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[68]
port 495 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 la_data_out[69]
port 496 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[6]
port 497 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[70]
port 498 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[71]
port 499 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 la_data_out[72]
port 500 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[73]
port 501 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[74]
port 502 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[75]
port 503 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[76]
port 504 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[77]
port 505 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[78]
port 506 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[79]
port 507 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 la_data_out[7]
port 508 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 la_data_out[80]
port 509 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[81]
port 510 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[82]
port 511 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[83]
port 512 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[84]
port 513 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[85]
port 514 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[86]
port 515 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[87]
port 516 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[88]
port 517 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[89]
port 518 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[8]
port 519 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[90]
port 520 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[91]
port 521 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 la_data_out[92]
port 522 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[93]
port 523 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[94]
port 524 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[95]
port 525 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 la_data_out[96]
port 526 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 la_data_out[97]
port 527 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[98]
port 528 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[99]
port 529 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la_data_out[9]
port 530 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 la_oenb[0]
port 531 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_oenb[100]
port 532 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[101]
port 533 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[102]
port 534 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[103]
port 535 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[104]
port 536 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oenb[105]
port 537 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[106]
port 538 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oenb[107]
port 539 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[108]
port 540 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[109]
port 541 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[10]
port 542 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[110]
port 543 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[111]
port 544 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[112]
port 545 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[113]
port 546 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_oenb[114]
port 547 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_oenb[115]
port 548 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[116]
port 549 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_oenb[117]
port 550 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[118]
port 551 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[119]
port 552 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[11]
port 553 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[120]
port 554 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_oenb[121]
port 555 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_oenb[122]
port 556 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[123]
port 557 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[124]
port 558 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_oenb[125]
port 559 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_oenb[126]
port 560 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oenb[127]
port 561 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[12]
port 562 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[13]
port 563 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[14]
port 564 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[15]
port 565 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[16]
port 566 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_oenb[17]
port 567 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[18]
port 568 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[19]
port 569 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[1]
port 570 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[20]
port 571 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[21]
port 572 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[22]
port 573 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[23]
port 574 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_oenb[24]
port 575 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[25]
port 576 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_oenb[26]
port 577 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[27]
port 578 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[28]
port 579 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[29]
port 580 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[2]
port 581 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[30]
port 582 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[31]
port 583 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[32]
port 584 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_oenb[33]
port 585 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_oenb[34]
port 586 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[35]
port 587 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_oenb[36]
port 588 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[37]
port 589 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[38]
port 590 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[39]
port 591 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[3]
port 592 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[40]
port 593 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[41]
port 594 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_oenb[42]
port 595 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_oenb[43]
port 596 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[44]
port 597 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_oenb[45]
port 598 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[46]
port 599 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[47]
port 600 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_oenb[48]
port 601 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[49]
port 602 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_oenb[4]
port 603 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_oenb[50]
port 604 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_oenb[51]
port 605 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_oenb[52]
port 606 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[53]
port 607 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[54]
port 608 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[55]
port 609 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[56]
port 610 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[57]
port 611 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_oenb[58]
port 612 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[59]
port 613 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_oenb[5]
port 614 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_oenb[60]
port 615 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[61]
port 616 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oenb[62]
port 617 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[63]
port 618 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[64]
port 619 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[65]
port 620 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[66]
port 621 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[67]
port 622 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[68]
port 623 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_oenb[69]
port 624 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_oenb[6]
port 625 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[70]
port 626 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[71]
port 627 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_oenb[72]
port 628 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oenb[73]
port 629 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[74]
port 630 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_oenb[75]
port 631 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[76]
port 632 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[77]
port 633 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[78]
port 634 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[79]
port 635 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[7]
port 636 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[80]
port 637 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[81]
port 638 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[82]
port 639 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[83]
port 640 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[84]
port 641 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[85]
port 642 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[86]
port 643 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[87]
port 644 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[88]
port 645 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_oenb[89]
port 646 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[8]
port 647 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[90]
port 648 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[91]
port 649 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[92]
port 650 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[93]
port 651 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[94]
port 652 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[95]
port 653 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_oenb[96]
port 654 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_oenb[97]
port 655 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_oenb[98]
port 656 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oenb[99]
port 657 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[9]
port 658 nsew signal input
rlabel metal2 s 118238 121102 118294 121902 6 user_irq[0]
port 659 nsew signal output
rlabel metal2 s 118790 121102 118846 121902 6 user_irq[1]
port 660 nsew signal output
rlabel metal2 s 119434 121102 119490 121902 6 user_irq[2]
port 661 nsew signal output
rlabel metal4 s 4208 2128 4528 119728 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 119728 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 119728 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 119728 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 119728 6 vssd1
port 663 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 119728 6 vssd1
port 663 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 119728 6 vssd1
port 663 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 119728 6 vssd1
port 663 nsew ground bidirectional
rlabel metal2 s 18 0 74 800 6 wb_clk_i
port 664 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_rst_i
port 665 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_uart_ack
port 666 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_uart_adr[0]
port 667 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wb_uart_adr[10]
port 668 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wb_uart_adr[11]
port 669 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wb_uart_adr[12]
port 670 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wb_uart_adr[13]
port 671 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wb_uart_adr[14]
port 672 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 wb_uart_adr[15]
port 673 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wb_uart_adr[16]
port 674 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wb_uart_adr[17]
port 675 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wb_uart_adr[18]
port 676 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wb_uart_adr[19]
port 677 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 wb_uart_adr[1]
port 678 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 wb_uart_adr[20]
port 679 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wb_uart_adr[21]
port 680 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wb_uart_adr[22]
port 681 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wb_uart_adr[23]
port 682 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wb_uart_adr[24]
port 683 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wb_uart_adr[25]
port 684 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wb_uart_adr[26]
port 685 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wb_uart_adr[27]
port 686 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wb_uart_adr[28]
port 687 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wb_uart_adr[29]
port 688 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wb_uart_adr[2]
port 689 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wb_uart_adr[30]
port 690 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wb_uart_adr[31]
port 691 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wb_uart_adr[3]
port 692 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 wb_uart_adr[4]
port 693 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 wb_uart_adr[5]
port 694 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wb_uart_adr[6]
port 695 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wb_uart_adr[7]
port 696 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 wb_uart_adr[8]
port 697 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wb_uart_adr[9]
port 698 nsew signal output
rlabel metal2 s 478 0 534 800 6 wb_uart_clk
port 699 nsew signal output
rlabel metal2 s 662 0 718 800 6 wb_uart_cyc
port 700 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 wb_uart_dat_fromcpu[0]
port 701 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wb_uart_dat_fromcpu[10]
port 702 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wb_uart_dat_fromcpu[11]
port 703 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wb_uart_dat_fromcpu[12]
port 704 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wb_uart_dat_fromcpu[13]
port 705 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wb_uart_dat_fromcpu[14]
port 706 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 wb_uart_dat_fromcpu[15]
port 707 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wb_uart_dat_fromcpu[16]
port 708 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 wb_uart_dat_fromcpu[17]
port 709 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wb_uart_dat_fromcpu[18]
port 710 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wb_uart_dat_fromcpu[19]
port 711 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 wb_uart_dat_fromcpu[1]
port 712 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wb_uart_dat_fromcpu[20]
port 713 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wb_uart_dat_fromcpu[21]
port 714 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wb_uart_dat_fromcpu[22]
port 715 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wb_uart_dat_fromcpu[23]
port 716 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 wb_uart_dat_fromcpu[24]
port 717 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wb_uart_dat_fromcpu[25]
port 718 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wb_uart_dat_fromcpu[26]
port 719 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wb_uart_dat_fromcpu[27]
port 720 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wb_uart_dat_fromcpu[28]
port 721 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wb_uart_dat_fromcpu[29]
port 722 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wb_uart_dat_fromcpu[2]
port 723 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 wb_uart_dat_fromcpu[30]
port 724 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wb_uart_dat_fromcpu[31]
port 725 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 wb_uart_dat_fromcpu[3]
port 726 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wb_uart_dat_fromcpu[4]
port 727 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wb_uart_dat_fromcpu[5]
port 728 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 wb_uart_dat_fromcpu[6]
port 729 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wb_uart_dat_fromcpu[7]
port 730 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wb_uart_dat_fromcpu[8]
port 731 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wb_uart_dat_fromcpu[9]
port 732 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 wb_uart_dat_tocpu[0]
port 733 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wb_uart_dat_tocpu[10]
port 734 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wb_uart_dat_tocpu[11]
port 735 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wb_uart_dat_tocpu[12]
port 736 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wb_uart_dat_tocpu[13]
port 737 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wb_uart_dat_tocpu[14]
port 738 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wb_uart_dat_tocpu[15]
port 739 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wb_uart_dat_tocpu[16]
port 740 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wb_uart_dat_tocpu[17]
port 741 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wb_uart_dat_tocpu[18]
port 742 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wb_uart_dat_tocpu[19]
port 743 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wb_uart_dat_tocpu[1]
port 744 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wb_uart_dat_tocpu[20]
port 745 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wb_uart_dat_tocpu[21]
port 746 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wb_uart_dat_tocpu[22]
port 747 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wb_uart_dat_tocpu[23]
port 748 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wb_uart_dat_tocpu[24]
port 749 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wb_uart_dat_tocpu[25]
port 750 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wb_uart_dat_tocpu[26]
port 751 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wb_uart_dat_tocpu[27]
port 752 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wb_uart_dat_tocpu[28]
port 753 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wb_uart_dat_tocpu[29]
port 754 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wb_uart_dat_tocpu[2]
port 755 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wb_uart_dat_tocpu[30]
port 756 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wb_uart_dat_tocpu[31]
port 757 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wb_uart_dat_tocpu[3]
port 758 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wb_uart_dat_tocpu[4]
port 759 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wb_uart_dat_tocpu[5]
port 760 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wb_uart_dat_tocpu[6]
port 761 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wb_uart_dat_tocpu[7]
port 762 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wb_uart_dat_tocpu[8]
port 763 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wb_uart_dat_tocpu[9]
port 764 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_uart_rst
port 765 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 wb_uart_sel[0]
port 766 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wb_uart_sel[1]
port 767 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wb_uart_sel[2]
port 768 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 wb_uart_sel[3]
port 769 nsew signal output
rlabel metal2 s 1030 0 1086 800 6 wb_uart_stb
port 770 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wb_uart_we
port 771 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_ack_o
port 772 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[0]
port 773 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[10]
port 774 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[11]
port 775 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_adr_i[12]
port 776 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[13]
port 777 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[14]
port 778 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[15]
port 779 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[16]
port 780 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[17]
port 781 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[18]
port 782 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[19]
port 783 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[1]
port 784 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[20]
port 785 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_adr_i[21]
port 786 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[22]
port 787 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[23]
port 788 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[24]
port 789 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_adr_i[25]
port 790 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[26]
port 791 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[27]
port 792 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[28]
port 793 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[29]
port 794 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[2]
port 795 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_adr_i[30]
port 796 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[31]
port 797 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[3]
port 798 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[4]
port 799 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_adr_i[5]
port 800 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[6]
port 801 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[7]
port 802 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[8]
port 803 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[9]
port 804 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_cyc_i
port 805 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[0]
port 806 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[10]
port 807 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[11]
port 808 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_i[12]
port 809 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_i[13]
port 810 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[14]
port 811 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[15]
port 812 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[16]
port 813 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[17]
port 814 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[18]
port 815 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[19]
port 816 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_i[1]
port 817 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_i[20]
port 818 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[21]
port 819 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[22]
port 820 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_i[23]
port 821 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[24]
port 822 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[25]
port 823 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_i[26]
port 824 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_i[27]
port 825 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_i[28]
port 826 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[29]
port 827 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[2]
port 828 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[30]
port 829 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[31]
port 830 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[3]
port 831 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[4]
port 832 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[5]
port 833 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[6]
port 834 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[7]
port 835 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[8]
port 836 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[9]
port 837 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[0]
port 838 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[10]
port 839 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[11]
port 840 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_o[12]
port 841 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[13]
port 842 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[14]
port 843 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_o[15]
port 844 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[16]
port 845 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_o[17]
port 846 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[18]
port 847 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_o[19]
port 848 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[1]
port 849 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[20]
port 850 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[21]
port 851 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_o[22]
port 852 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[23]
port 853 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[24]
port 854 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[25]
port 855 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_o[26]
port 856 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[27]
port 857 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_o[28]
port 858 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_o[29]
port 859 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[2]
port 860 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[30]
port 861 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_o[31]
port 862 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[3]
port 863 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[4]
port 864 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[5]
port 865 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[6]
port 866 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_o[7]
port 867 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[8]
port 868 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[9]
port 869 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_sel_i[0]
port 870 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_sel_i[1]
port 871 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_sel_i[2]
port 872 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_sel_i[3]
port 873 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_stb_i
port 874 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_we_i
port 875 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 119758 121902
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 38817546
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc/openlane/rvj1_caravel_soc/runs/rvj1_caravel_soc/results/signoff/rvj1_caravel_soc.magic.gds
string GDS_START 1262256
<< end >>

