VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rvj1_caravel_soc
  CLASS BLOCK ;
  FOREIGN rvj1_caravel_soc ;
  ORIGIN 0.000 0.000 ;
  SIZE 591.480 BY 602.200 ;
  PIN dram_addr0[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END dram_addr0[-1]
  PIN dram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 183.640 591.480 184.240 ;
    END
  END dram_addr0[0]
  PIN dram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 299.240 591.480 299.840 ;
    END
  END dram_clk0
  PIN dram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 421.640 591.480 422.240 ;
    END
  END dram_csb0
  PIN dram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 20.440 591.480 21.040 ;
    END
  END dram_din0[0]
  PIN dram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 598.200 480.150 602.200 ;
    END
  END dram_din0[10]
  PIN dram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 598.200 332.030 602.200 ;
    END
  END dram_din0[11]
  PIN dram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END dram_din0[12]
  PIN dram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 380.840 591.480 381.440 ;
    END
  END dram_din0[13]
  PIN dram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 598.200 383.550 602.200 ;
    END
  END dram_din0[14]
  PIN dram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 598.200 364.230 602.200 ;
    END
  END dram_din0[15]
  PIN dram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END dram_din0[16]
  PIN dram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END dram_din0[17]
  PIN dram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 115.640 591.480 116.240 ;
    END
  END dram_din0[18]
  PIN dram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END dram_din0[19]
  PIN dram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 292.440 591.480 293.040 ;
    END
  END dram_din0[1]
  PIN dram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 598.200 299.830 602.200 ;
    END
  END dram_din0[20]
  PIN dram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 61.240 591.480 61.840 ;
    END
  END dram_din0[21]
  PIN dram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END dram_din0[22]
  PIN dram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END dram_din0[23]
  PIN dram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END dram_din0[24]
  PIN dram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 428.440 591.480 429.040 ;
    END
  END dram_din0[25]
  PIN dram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END dram_din0[26]
  PIN dram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 74.840 591.480 75.440 ;
    END
  END dram_din0[27]
  PIN dram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 598.200 435.070 602.200 ;
    END
  END dram_din0[28]
  PIN dram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 598.200 563.870 602.200 ;
    END
  END dram_din0[29]
  PIN dram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 448.840 591.480 449.440 ;
    END
  END dram_din0[2]
  PIN dram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 598.200 48.670 602.200 ;
    END
  END dram_din0[30]
  PIN dram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END dram_din0[31]
  PIN dram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 13.640 591.480 14.240 ;
    END
  END dram_din0[3]
  PIN dram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 244.840 591.480 245.440 ;
    END
  END dram_din0[4]
  PIN dram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END dram_din0[5]
  PIN dram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END dram_din0[6]
  PIN dram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END dram_din0[7]
  PIN dram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END dram_din0[8]
  PIN dram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 598.200 106.630 602.200 ;
    END
  END dram_din0[9]
  PIN dram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 598.200 100.190 602.200 ;
    END
  END dram_dout0[0]
  PIN dram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END dram_dout0[10]
  PIN dram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END dram_dout0[11]
  PIN dram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 503.240 591.480 503.840 ;
    END
  END dram_dout0[12]
  PIN dram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 40.840 591.480 41.440 ;
    END
  END dram_dout0[13]
  PIN dram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 265.240 591.480 265.840 ;
    END
  END dram_dout0[14]
  PIN dram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END dram_dout0[15]
  PIN dram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END dram_dout0[16]
  PIN dram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 598.200 525.230 602.200 ;
    END
  END dram_dout0[17]
  PIN dram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END dram_dout0[18]
  PIN dram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 598.200 357.790 602.200 ;
    END
  END dram_dout0[19]
  PIN dram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 149.640 591.480 150.240 ;
    END
  END dram_dout0[1]
  PIN dram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END dram_dout0[20]
  PIN dram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 251.640 591.480 252.240 ;
    END
  END dram_dout0[21]
  PIN dram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END dram_dout0[22]
  PIN dram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END dram_dout0[23]
  PIN dram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 598.200 538.110 602.200 ;
    END
  END dram_dout0[24]
  PIN dram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 598.200 235.430 602.200 ;
    END
  END dram_dout0[25]
  PIN dram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END dram_dout0[26]
  PIN dram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END dram_dout0[27]
  PIN dram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END dram_dout0[28]
  PIN dram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 258.440 591.480 259.040 ;
    END
  END dram_dout0[29]
  PIN dram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END dram_dout0[2]
  PIN dram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END dram_dout0[30]
  PIN dram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 598.200 216.110 602.200 ;
    END
  END dram_dout0[31]
  PIN dram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 469.240 591.480 469.840 ;
    END
  END dram_dout0[3]
  PIN dram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END dram_dout0[4]
  PIN dram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 598.200 370.670 602.200 ;
    END
  END dram_dout0[5]
  PIN dram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END dram_dout0[6]
  PIN dram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END dram_dout0[7]
  PIN dram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 197.240 591.480 197.840 ;
    END
  END dram_dout0[8]
  PIN dram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END dram_dout0[9]
  PIN dram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 489.640 591.480 490.240 ;
    END
  END dram_web0
  PIN dram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END dram_wmask0[0]
  PIN dram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 598.200 409.310 602.200 ;
    END
  END dram_wmask0[1]
  PIN dram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END dram_wmask0[2]
  PIN dram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END dram_wmask0[3]
  PIN iram_addr0[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END iram_addr0[-1]
  PIN iram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 598.200 151.710 602.200 ;
    END
  END iram_addr0[0]
  PIN iram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 408.040 591.480 408.640 ;
    END
  END iram_clk0
  PIN iram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END iram_csb0
  PIN iram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 598.200 402.870 602.200 ;
    END
  END iram_din0[0]
  PIN iram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 102.040 591.480 102.640 ;
    END
  END iram_din0[10]
  PIN iram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END iram_din0[11]
  PIN iram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END iram_din0[12]
  PIN iram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 367.240 591.480 367.840 ;
    END
  END iram_din0[13]
  PIN iram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END iram_din0[14]
  PIN iram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 136.040 591.480 136.640 ;
    END
  END iram_din0[15]
  PIN iram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END iram_din0[16]
  PIN iram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 374.040 591.480 374.640 ;
    END
  END iram_din0[17]
  PIN iram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 598.200 171.030 602.200 ;
    END
  END iram_din0[18]
  PIN iram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END iram_din0[19]
  PIN iram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END iram_din0[1]
  PIN iram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 598.200 55.110 602.200 ;
    END
  END iram_din0[20]
  PIN iram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 598.200 428.630 602.200 ;
    END
  END iram_din0[21]
  PIN iram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END iram_din0[22]
  PIN iram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 401.240 591.480 401.840 ;
    END
  END iram_din0[23]
  PIN iram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END iram_din0[24]
  PIN iram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END iram_din0[25]
  PIN iram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END iram_din0[26]
  PIN iram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 598.200 293.390 602.200 ;
    END
  END iram_din0[27]
  PIN iram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 571.240 591.480 571.840 ;
    END
  END iram_din0[28]
  PIN iram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END iram_din0[29]
  PIN iram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 163.240 591.480 163.840 ;
    END
  END iram_din0[2]
  PIN iram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END iram_din0[30]
  PIN iram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 598.200 274.070 602.200 ;
    END
  END iram_din0[31]
  PIN iram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 598.200 312.710 602.200 ;
    END
  END iram_din0[3]
  PIN iram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 204.040 591.480 204.640 ;
    END
  END iram_din0[4]
  PIN iram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 346.840 591.480 347.440 ;
    END
  END iram_din0[5]
  PIN iram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END iram_din0[6]
  PIN iram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END iram_din0[7]
  PIN iram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 598.200 486.590 602.200 ;
    END
  END iram_din0[8]
  PIN iram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END iram_din0[9]
  PIN iram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END iram_dout0[0]
  PIN iram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 476.040 591.480 476.640 ;
    END
  END iram_dout0[10]
  PIN iram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END iram_dout0[11]
  PIN iram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END iram_dout0[12]
  PIN iram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 598.200 505.910 602.200 ;
    END
  END iram_dout0[13]
  PIN iram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 81.640 591.480 82.240 ;
    END
  END iram_dout0[14]
  PIN iram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END iram_dout0[15]
  PIN iram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END iram_dout0[16]
  PIN iram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 88.440 591.480 89.040 ;
    END
  END iram_dout0[17]
  PIN iram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END iram_dout0[18]
  PIN iram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 598.200 42.230 602.200 ;
    END
  END iram_dout0[19]
  PIN iram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END iram_dout0[1]
  PIN iram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 598.200 261.190 602.200 ;
    END
  END iram_dout0[20]
  PIN iram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 564.440 591.480 565.040 ;
    END
  END iram_dout0[21]
  PIN iram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 360.440 591.480 361.040 ;
    END
  END iram_dout0[22]
  PIN iram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END iram_dout0[23]
  PIN iram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 598.200 454.390 602.200 ;
    END
  END iram_dout0[24]
  PIN iram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END iram_dout0[25]
  PIN iram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 598.200 138.830 602.200 ;
    END
  END iram_dout0[26]
  PIN iram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END iram_dout0[27]
  PIN iram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 598.200 35.790 602.200 ;
    END
  END iram_dout0[28]
  PIN iram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END iram_dout0[29]
  PIN iram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 598.200 473.710 602.200 ;
    END
  END iram_dout0[2]
  PIN iram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END iram_dout0[30]
  PIN iram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 108.840 591.480 109.440 ;
    END
  END iram_dout0[31]
  PIN iram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END iram_dout0[3]
  PIN iram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 598.200 377.110 602.200 ;
    END
  END iram_dout0[4]
  PIN iram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 190.440 591.480 191.040 ;
    END
  END iram_dout0[5]
  PIN iram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END iram_dout0[6]
  PIN iram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 27.240 591.480 27.840 ;
    END
  END iram_dout0[7]
  PIN iram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 598.200 93.750 602.200 ;
    END
  END iram_dout0[8]
  PIN iram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END iram_dout0[9]
  PIN iram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END iram_web0
  PIN iram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END iram_wmask0[0]
  PIN iram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 598.200 415.750 602.200 ;
    END
  END iram_wmask0[1]
  PIN iram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END iram_wmask0[2]
  PIN iram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 598.200 550.990 602.200 ;
    END
  END iram_wmask0[3]
  PIN jedro_1_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END jedro_1_rstn
  PIN sel_wb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END sel_wb
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 590.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 590.480 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 598.200 254.750 602.200 ;
    END
  END wb_rst_i
  PIN wb_uart_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 591.640 591.480 592.240 ;
    END
  END wb_uart_ack
  PIN wb_uart_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 598.200 544.550 602.200 ;
    END
  END wb_uart_adr[0]
  PIN wb_uart_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END wb_uart_adr[10]
  PIN wb_uart_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 598.200 196.790 602.200 ;
    END
  END wb_uart_adr[11]
  PIN wb_uart_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 510.040 591.480 510.640 ;
    END
  END wb_uart_adr[12]
  PIN wb_uart_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 598.200 10.030 602.200 ;
    END
  END wb_uart_adr[13]
  PIN wb_uart_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END wb_uart_adr[14]
  PIN wb_uart_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 598.200 113.070 602.200 ;
    END
  END wb_uart_adr[15]
  PIN wb_uart_adr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END wb_uart_adr[16]
  PIN wb_uart_adr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wb_uart_adr[17]
  PIN wb_uart_adr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 598.200 119.510 602.200 ;
    END
  END wb_uart_adr[18]
  PIN wb_uart_adr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wb_uart_adr[19]
  PIN wb_uart_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 598.200 512.350 602.200 ;
    END
  END wb_uart_adr[1]
  PIN wb_uart_adr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END wb_uart_adr[20]
  PIN wb_uart_adr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END wb_uart_adr[21]
  PIN wb_uart_adr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 598.200 3.590 602.200 ;
    END
  END wb_uart_adr[22]
  PIN wb_uart_adr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 598.200 557.430 602.200 ;
    END
  END wb_uart_adr[23]
  PIN wb_uart_adr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END wb_uart_adr[24]
  PIN wb_uart_adr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wb_uart_adr[25]
  PIN wb_uart_adr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wb_uart_adr[26]
  PIN wb_uart_adr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 598.200 351.350 602.200 ;
    END
  END wb_uart_adr[27]
  PIN wb_uart_adr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 598.200 447.950 602.200 ;
    END
  END wb_uart_adr[28]
  PIN wb_uart_adr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wb_uart_adr[29]
  PIN wb_uart_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 34.040 591.480 34.640 ;
    END
  END wb_uart_adr[2]
  PIN wb_uart_adr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 578.040 591.480 578.640 ;
    END
  END wb_uart_adr[30]
  PIN wb_uart_adr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END wb_uart_adr[31]
  PIN wb_uart_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wb_uart_adr[3]
  PIN wb_uart_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 231.240 591.480 231.840 ;
    END
  END wb_uart_adr[4]
  PIN wb_uart_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 550.840 591.480 551.440 ;
    END
  END wb_uart_adr[5]
  PIN wb_uart_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 598.200 158.150 602.200 ;
    END
  END wb_uart_adr[6]
  PIN wb_uart_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END wb_uart_adr[7]
  PIN wb_uart_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END wb_uart_adr[8]
  PIN wb_uart_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 68.040 591.480 68.640 ;
    END
  END wb_uart_adr[9]
  PIN wb_uart_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END wb_uart_clk
  PIN wb_uart_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END wb_uart_cyc
  PIN wb_uart_dat_fromcpu[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 176.840 591.480 177.440 ;
    END
  END wb_uart_dat_fromcpu[0]
  PIN wb_uart_dat_fromcpu[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 122.440 591.480 123.040 ;
    END
  END wb_uart_dat_fromcpu[10]
  PIN wb_uart_dat_fromcpu[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 598.200 80.870 602.200 ;
    END
  END wb_uart_dat_fromcpu[11]
  PIN wb_uart_dat_fromcpu[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wb_uart_dat_fromcpu[12]
  PIN wb_uart_dat_fromcpu[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END wb_uart_dat_fromcpu[13]
  PIN wb_uart_dat_fromcpu[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 598.200 228.990 602.200 ;
    END
  END wb_uart_dat_fromcpu[14]
  PIN wb_uart_dat_fromcpu[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END wb_uart_dat_fromcpu[15]
  PIN wb_uart_dat_fromcpu[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END wb_uart_dat_fromcpu[16]
  PIN wb_uart_dat_fromcpu[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wb_uart_dat_fromcpu[17]
  PIN wb_uart_dat_fromcpu[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wb_uart_dat_fromcpu[18]
  PIN wb_uart_dat_fromcpu[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 598.200 222.550 602.200 ;
    END
  END wb_uart_dat_fromcpu[19]
  PIN wb_uart_dat_fromcpu[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END wb_uart_dat_fromcpu[1]
  PIN wb_uart_dat_fromcpu[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 210.840 591.480 211.440 ;
    END
  END wb_uart_dat_fromcpu[20]
  PIN wb_uart_dat_fromcpu[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wb_uart_dat_fromcpu[21]
  PIN wb_uart_dat_fromcpu[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 544.040 591.480 544.640 ;
    END
  END wb_uart_dat_fromcpu[22]
  PIN wb_uart_dat_fromcpu[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 598.200 570.310 602.200 ;
    END
  END wb_uart_dat_fromcpu[23]
  PIN wb_uart_dat_fromcpu[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wb_uart_dat_fromcpu[24]
  PIN wb_uart_dat_fromcpu[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 272.040 591.480 272.640 ;
    END
  END wb_uart_dat_fromcpu[25]
  PIN wb_uart_dat_fromcpu[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END wb_uart_dat_fromcpu[26]
  PIN wb_uart_dat_fromcpu[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 598.200 531.670 602.200 ;
    END
  END wb_uart_dat_fromcpu[27]
  PIN wb_uart_dat_fromcpu[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wb_uart_dat_fromcpu[28]
  PIN wb_uart_dat_fromcpu[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 224.440 591.480 225.040 ;
    END
  END wb_uart_dat_fromcpu[29]
  PIN wb_uart_dat_fromcpu[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 462.440 591.480 463.040 ;
    END
  END wb_uart_dat_fromcpu[2]
  PIN wb_uart_dat_fromcpu[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 496.440 591.480 497.040 ;
    END
  END wb_uart_dat_fromcpu[30]
  PIN wb_uart_dat_fromcpu[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 414.840 591.480 415.440 ;
    END
  END wb_uart_dat_fromcpu[31]
  PIN wb_uart_dat_fromcpu[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 598.200 132.390 602.200 ;
    END
  END wb_uart_dat_fromcpu[3]
  PIN wb_uart_dat_fromcpu[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 598.200 61.550 602.200 ;
    END
  END wb_uart_dat_fromcpu[4]
  PIN wb_uart_dat_fromcpu[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END wb_uart_dat_fromcpu[5]
  PIN wb_uart_dat_fromcpu[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 557.640 591.480 558.240 ;
    END
  END wb_uart_dat_fromcpu[6]
  PIN wb_uart_dat_fromcpu[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 598.200 319.150 602.200 ;
    END
  END wb_uart_dat_fromcpu[7]
  PIN wb_uart_dat_fromcpu[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wb_uart_dat_fromcpu[8]
  PIN wb_uart_dat_fromcpu[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 598.200 280.510 602.200 ;
    END
  END wb_uart_dat_fromcpu[9]
  PIN wb_uart_dat_tocpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wb_uart_dat_tocpu[0]
  PIN wb_uart_dat_tocpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END wb_uart_dat_tocpu[10]
  PIN wb_uart_dat_tocpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 523.640 591.480 524.240 ;
    END
  END wb_uart_dat_tocpu[11]
  PIN wb_uart_dat_tocpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 598.200 209.670 602.200 ;
    END
  END wb_uart_dat_tocpu[12]
  PIN wb_uart_dat_tocpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 598.200 338.470 602.200 ;
    END
  END wb_uart_dat_tocpu[13]
  PIN wb_uart_dat_tocpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END wb_uart_dat_tocpu[14]
  PIN wb_uart_dat_tocpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wb_uart_dat_tocpu[15]
  PIN wb_uart_dat_tocpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wb_uart_dat_tocpu[16]
  PIN wb_uart_dat_tocpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 598.200 583.190 602.200 ;
    END
  END wb_uart_dat_tocpu[17]
  PIN wb_uart_dat_tocpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END wb_uart_dat_tocpu[18]
  PIN wb_uart_dat_tocpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wb_uart_dat_tocpu[19]
  PIN wb_uart_dat_tocpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END wb_uart_dat_tocpu[1]
  PIN wb_uart_dat_tocpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END wb_uart_dat_tocpu[20]
  PIN wb_uart_dat_tocpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 598.200 164.590 602.200 ;
    END
  END wb_uart_dat_tocpu[21]
  PIN wb_uart_dat_tocpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END wb_uart_dat_tocpu[22]
  PIN wb_uart_dat_tocpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 598.200 306.270 602.200 ;
    END
  END wb_uart_dat_tocpu[23]
  PIN wb_uart_dat_tocpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 598.200 29.350 602.200 ;
    END
  END wb_uart_dat_tocpu[24]
  PIN wb_uart_dat_tocpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END wb_uart_dat_tocpu[25]
  PIN wb_uart_dat_tocpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END wb_uart_dat_tocpu[26]
  PIN wb_uart_dat_tocpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 598.200 177.470 602.200 ;
    END
  END wb_uart_dat_tocpu[27]
  PIN wb_uart_dat_tocpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END wb_uart_dat_tocpu[28]
  PIN wb_uart_dat_tocpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 598.200 16.470 602.200 ;
    END
  END wb_uart_dat_tocpu[29]
  PIN wb_uart_dat_tocpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END wb_uart_dat_tocpu[2]
  PIN wb_uart_dat_tocpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 598.200 22.910 602.200 ;
    END
  END wb_uart_dat_tocpu[30]
  PIN wb_uart_dat_tocpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END wb_uart_dat_tocpu[31]
  PIN wb_uart_dat_tocpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 598.200 248.310 602.200 ;
    END
  END wb_uart_dat_tocpu[3]
  PIN wb_uart_dat_tocpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wb_uart_dat_tocpu[4]
  PIN wb_uart_dat_tocpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END wb_uart_dat_tocpu[5]
  PIN wb_uart_dat_tocpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 598.200 67.990 602.200 ;
    END
  END wb_uart_dat_tocpu[6]
  PIN wb_uart_dat_tocpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 326.440 591.480 327.040 ;
    END
  END wb_uart_dat_tocpu[7]
  PIN wb_uart_dat_tocpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wb_uart_dat_tocpu[8]
  PIN wb_uart_dat_tocpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END wb_uart_dat_tocpu[9]
  PIN wb_uart_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END wb_uart_rst
  PIN wb_uart_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wb_uart_sel[0]
  PIN wb_uart_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 394.440 591.480 395.040 ;
    END
  END wb_uart_sel[1]
  PIN wb_uart_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END wb_uart_sel[2]
  PIN wb_uart_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 598.200 286.950 602.200 ;
    END
  END wb_uart_sel[3]
  PIN wb_uart_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 54.440 591.480 55.040 ;
    END
  END wb_uart_stb
  PIN wb_uart_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 598.200 203.230 602.200 ;
    END
  END wb_uart_we
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 598.200 467.270 602.200 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 598.200 344.910 602.200 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 598.200 125.950 602.200 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 387.640 591.480 388.240 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 353.640 591.480 354.240 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 312.840 591.480 313.440 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 142.840 591.480 143.440 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 584.840 591.480 585.440 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 95.240 591.480 95.840 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 598.200 145.270 602.200 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 598.200 267.630 602.200 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 306.040 591.480 306.640 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 530.440 591.480 531.040 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 217.640 591.480 218.240 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 598.200 499.470 602.200 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 129.240 591.480 129.840 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 598.200 241.870 602.200 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 482.840 591.480 483.440 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 278.840 591.480 279.440 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 598.200 576.750 602.200 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 598.200 87.310 602.200 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 333.240 591.480 333.840 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 598.200 589.630 602.200 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 442.040 591.480 442.640 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 170.040 591.480 170.640 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 598.200 518.790 602.200 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 340.040 591.480 340.640 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 0.040 591.480 0.640 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 238.040 591.480 238.640 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 598.200 493.030 602.200 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 516.840 591.480 517.440 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 6.840 591.480 7.440 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 319.640 591.480 320.240 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 537.240 591.480 537.840 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 598.200 460.830 602.200 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 47.640 591.480 48.240 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 598.200 441.510 602.200 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 598.200 183.910 602.200 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 598.200 325.590 602.200 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 598.200 190.350 602.200 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 598.200 422.190 602.200 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 156.440 591.480 157.040 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 455.640 591.480 456.240 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 435.240 591.480 435.840 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 598.200 396.430 602.200 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 598.200 389.990 602.200 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 598.200 74.430 602.200 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 285.640 591.480 286.240 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 585.580 590.325 ;
      LAYER met1 ;
        RECT 0.070 4.460 591.030 595.640 ;
      LAYER met2 ;
        RECT 0.100 597.920 3.030 600.965 ;
        RECT 3.870 597.920 9.470 600.965 ;
        RECT 10.310 597.920 15.910 600.965 ;
        RECT 16.750 597.920 22.350 600.965 ;
        RECT 23.190 597.920 28.790 600.965 ;
        RECT 29.630 597.920 35.230 600.965 ;
        RECT 36.070 597.920 41.670 600.965 ;
        RECT 42.510 597.920 48.110 600.965 ;
        RECT 48.950 597.920 54.550 600.965 ;
        RECT 55.390 597.920 60.990 600.965 ;
        RECT 61.830 597.920 67.430 600.965 ;
        RECT 68.270 597.920 73.870 600.965 ;
        RECT 74.710 597.920 80.310 600.965 ;
        RECT 81.150 597.920 86.750 600.965 ;
        RECT 87.590 597.920 93.190 600.965 ;
        RECT 94.030 597.920 99.630 600.965 ;
        RECT 100.470 597.920 106.070 600.965 ;
        RECT 106.910 597.920 112.510 600.965 ;
        RECT 113.350 597.920 118.950 600.965 ;
        RECT 119.790 597.920 125.390 600.965 ;
        RECT 126.230 597.920 131.830 600.965 ;
        RECT 132.670 597.920 138.270 600.965 ;
        RECT 139.110 597.920 144.710 600.965 ;
        RECT 145.550 597.920 151.150 600.965 ;
        RECT 151.990 597.920 157.590 600.965 ;
        RECT 158.430 597.920 164.030 600.965 ;
        RECT 164.870 597.920 170.470 600.965 ;
        RECT 171.310 597.920 176.910 600.965 ;
        RECT 177.750 597.920 183.350 600.965 ;
        RECT 184.190 597.920 189.790 600.965 ;
        RECT 190.630 597.920 196.230 600.965 ;
        RECT 197.070 597.920 202.670 600.965 ;
        RECT 203.510 597.920 209.110 600.965 ;
        RECT 209.950 597.920 215.550 600.965 ;
        RECT 216.390 597.920 221.990 600.965 ;
        RECT 222.830 597.920 228.430 600.965 ;
        RECT 229.270 597.920 234.870 600.965 ;
        RECT 235.710 597.920 241.310 600.965 ;
        RECT 242.150 597.920 247.750 600.965 ;
        RECT 248.590 597.920 254.190 600.965 ;
        RECT 255.030 597.920 260.630 600.965 ;
        RECT 261.470 597.920 267.070 600.965 ;
        RECT 267.910 597.920 273.510 600.965 ;
        RECT 274.350 597.920 279.950 600.965 ;
        RECT 280.790 597.920 286.390 600.965 ;
        RECT 287.230 597.920 292.830 600.965 ;
        RECT 293.670 597.920 299.270 600.965 ;
        RECT 300.110 597.920 305.710 600.965 ;
        RECT 306.550 597.920 312.150 600.965 ;
        RECT 312.990 597.920 318.590 600.965 ;
        RECT 319.430 597.920 325.030 600.965 ;
        RECT 325.870 597.920 331.470 600.965 ;
        RECT 332.310 597.920 337.910 600.965 ;
        RECT 338.750 597.920 344.350 600.965 ;
        RECT 345.190 597.920 350.790 600.965 ;
        RECT 351.630 597.920 357.230 600.965 ;
        RECT 358.070 597.920 363.670 600.965 ;
        RECT 364.510 597.920 370.110 600.965 ;
        RECT 370.950 597.920 376.550 600.965 ;
        RECT 377.390 597.920 382.990 600.965 ;
        RECT 383.830 597.920 389.430 600.965 ;
        RECT 390.270 597.920 395.870 600.965 ;
        RECT 396.710 597.920 402.310 600.965 ;
        RECT 403.150 597.920 408.750 600.965 ;
        RECT 409.590 597.920 415.190 600.965 ;
        RECT 416.030 597.920 421.630 600.965 ;
        RECT 422.470 597.920 428.070 600.965 ;
        RECT 428.910 597.920 434.510 600.965 ;
        RECT 435.350 597.920 440.950 600.965 ;
        RECT 441.790 597.920 447.390 600.965 ;
        RECT 448.230 597.920 453.830 600.965 ;
        RECT 454.670 597.920 460.270 600.965 ;
        RECT 461.110 597.920 466.710 600.965 ;
        RECT 467.550 597.920 473.150 600.965 ;
        RECT 473.990 597.920 479.590 600.965 ;
        RECT 480.430 597.920 486.030 600.965 ;
        RECT 486.870 597.920 492.470 600.965 ;
        RECT 493.310 597.920 498.910 600.965 ;
        RECT 499.750 597.920 505.350 600.965 ;
        RECT 506.190 597.920 511.790 600.965 ;
        RECT 512.630 597.920 518.230 600.965 ;
        RECT 519.070 597.920 524.670 600.965 ;
        RECT 525.510 597.920 531.110 600.965 ;
        RECT 531.950 597.920 537.550 600.965 ;
        RECT 538.390 597.920 543.990 600.965 ;
        RECT 544.830 597.920 550.430 600.965 ;
        RECT 551.270 597.920 556.870 600.965 ;
        RECT 557.710 597.920 563.310 600.965 ;
        RECT 564.150 597.920 569.750 600.965 ;
        RECT 570.590 597.920 576.190 600.965 ;
        RECT 577.030 597.920 582.630 600.965 ;
        RECT 583.470 597.920 589.070 600.965 ;
        RECT 589.910 597.920 591.000 600.965 ;
        RECT 0.100 4.280 591.000 597.920 ;
        RECT 0.650 0.155 6.250 4.280 ;
        RECT 7.090 0.155 12.690 4.280 ;
        RECT 13.530 0.155 19.130 4.280 ;
        RECT 19.970 0.155 25.570 4.280 ;
        RECT 26.410 0.155 32.010 4.280 ;
        RECT 32.850 0.155 38.450 4.280 ;
        RECT 39.290 0.155 44.890 4.280 ;
        RECT 45.730 0.155 51.330 4.280 ;
        RECT 52.170 0.155 57.770 4.280 ;
        RECT 58.610 0.155 64.210 4.280 ;
        RECT 65.050 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 83.530 4.280 ;
        RECT 84.370 0.155 89.970 4.280 ;
        RECT 90.810 0.155 96.410 4.280 ;
        RECT 97.250 0.155 102.850 4.280 ;
        RECT 103.690 0.155 109.290 4.280 ;
        RECT 110.130 0.155 115.730 4.280 ;
        RECT 116.570 0.155 122.170 4.280 ;
        RECT 123.010 0.155 128.610 4.280 ;
        RECT 129.450 0.155 135.050 4.280 ;
        RECT 135.890 0.155 141.490 4.280 ;
        RECT 142.330 0.155 147.930 4.280 ;
        RECT 148.770 0.155 154.370 4.280 ;
        RECT 155.210 0.155 160.810 4.280 ;
        RECT 161.650 0.155 167.250 4.280 ;
        RECT 168.090 0.155 173.690 4.280 ;
        RECT 174.530 0.155 180.130 4.280 ;
        RECT 180.970 0.155 186.570 4.280 ;
        RECT 187.410 0.155 193.010 4.280 ;
        RECT 193.850 0.155 199.450 4.280 ;
        RECT 200.290 0.155 205.890 4.280 ;
        RECT 206.730 0.155 212.330 4.280 ;
        RECT 213.170 0.155 218.770 4.280 ;
        RECT 219.610 0.155 225.210 4.280 ;
        RECT 226.050 0.155 231.650 4.280 ;
        RECT 232.490 0.155 238.090 4.280 ;
        RECT 238.930 0.155 244.530 4.280 ;
        RECT 245.370 0.155 250.970 4.280 ;
        RECT 251.810 0.155 257.410 4.280 ;
        RECT 258.250 0.155 263.850 4.280 ;
        RECT 264.690 0.155 270.290 4.280 ;
        RECT 271.130 0.155 276.730 4.280 ;
        RECT 277.570 0.155 283.170 4.280 ;
        RECT 284.010 0.155 289.610 4.280 ;
        RECT 290.450 0.155 296.050 4.280 ;
        RECT 296.890 0.155 302.490 4.280 ;
        RECT 303.330 0.155 308.930 4.280 ;
        RECT 309.770 0.155 315.370 4.280 ;
        RECT 316.210 0.155 321.810 4.280 ;
        RECT 322.650 0.155 328.250 4.280 ;
        RECT 329.090 0.155 334.690 4.280 ;
        RECT 335.530 0.155 341.130 4.280 ;
        RECT 341.970 0.155 347.570 4.280 ;
        RECT 348.410 0.155 354.010 4.280 ;
        RECT 354.850 0.155 360.450 4.280 ;
        RECT 361.290 0.155 366.890 4.280 ;
        RECT 367.730 0.155 373.330 4.280 ;
        RECT 374.170 0.155 379.770 4.280 ;
        RECT 380.610 0.155 386.210 4.280 ;
        RECT 387.050 0.155 392.650 4.280 ;
        RECT 393.490 0.155 399.090 4.280 ;
        RECT 399.930 0.155 405.530 4.280 ;
        RECT 406.370 0.155 411.970 4.280 ;
        RECT 412.810 0.155 418.410 4.280 ;
        RECT 419.250 0.155 424.850 4.280 ;
        RECT 425.690 0.155 431.290 4.280 ;
        RECT 432.130 0.155 437.730 4.280 ;
        RECT 438.570 0.155 444.170 4.280 ;
        RECT 445.010 0.155 450.610 4.280 ;
        RECT 451.450 0.155 457.050 4.280 ;
        RECT 457.890 0.155 463.490 4.280 ;
        RECT 464.330 0.155 469.930 4.280 ;
        RECT 470.770 0.155 476.370 4.280 ;
        RECT 477.210 0.155 482.810 4.280 ;
        RECT 483.650 0.155 489.250 4.280 ;
        RECT 490.090 0.155 495.690 4.280 ;
        RECT 496.530 0.155 502.130 4.280 ;
        RECT 502.970 0.155 508.570 4.280 ;
        RECT 509.410 0.155 515.010 4.280 ;
        RECT 515.850 0.155 521.450 4.280 ;
        RECT 522.290 0.155 527.890 4.280 ;
        RECT 528.730 0.155 534.330 4.280 ;
        RECT 535.170 0.155 540.770 4.280 ;
        RECT 541.610 0.155 547.210 4.280 ;
        RECT 548.050 0.155 553.650 4.280 ;
        RECT 554.490 0.155 560.090 4.280 ;
        RECT 560.930 0.155 566.530 4.280 ;
        RECT 567.370 0.155 572.970 4.280 ;
        RECT 573.810 0.155 579.410 4.280 ;
        RECT 580.250 0.155 585.850 4.280 ;
        RECT 586.690 0.155 591.000 4.280 ;
      LAYER met3 ;
        RECT 4.000 599.440 589.195 600.945 ;
        RECT 4.400 598.040 589.195 599.440 ;
        RECT 4.000 592.640 589.195 598.040 ;
        RECT 4.400 591.240 587.080 592.640 ;
        RECT 4.000 585.840 589.195 591.240 ;
        RECT 4.400 584.440 587.080 585.840 ;
        RECT 4.000 579.040 589.195 584.440 ;
        RECT 4.400 577.640 587.080 579.040 ;
        RECT 4.000 572.240 589.195 577.640 ;
        RECT 4.400 570.840 587.080 572.240 ;
        RECT 4.000 565.440 589.195 570.840 ;
        RECT 4.400 564.040 587.080 565.440 ;
        RECT 4.000 558.640 589.195 564.040 ;
        RECT 4.400 557.240 587.080 558.640 ;
        RECT 4.000 551.840 589.195 557.240 ;
        RECT 4.400 550.440 587.080 551.840 ;
        RECT 4.000 545.040 589.195 550.440 ;
        RECT 4.400 543.640 587.080 545.040 ;
        RECT 4.000 538.240 589.195 543.640 ;
        RECT 4.400 536.840 587.080 538.240 ;
        RECT 4.000 531.440 589.195 536.840 ;
        RECT 4.400 530.040 587.080 531.440 ;
        RECT 4.000 524.640 589.195 530.040 ;
        RECT 4.400 523.240 587.080 524.640 ;
        RECT 4.000 517.840 589.195 523.240 ;
        RECT 4.400 516.440 587.080 517.840 ;
        RECT 4.000 511.040 589.195 516.440 ;
        RECT 4.400 509.640 587.080 511.040 ;
        RECT 4.000 504.240 589.195 509.640 ;
        RECT 4.400 502.840 587.080 504.240 ;
        RECT 4.000 497.440 589.195 502.840 ;
        RECT 4.400 496.040 587.080 497.440 ;
        RECT 4.000 490.640 589.195 496.040 ;
        RECT 4.400 489.240 587.080 490.640 ;
        RECT 4.000 483.840 589.195 489.240 ;
        RECT 4.400 482.440 587.080 483.840 ;
        RECT 4.000 477.040 589.195 482.440 ;
        RECT 4.400 475.640 587.080 477.040 ;
        RECT 4.000 470.240 589.195 475.640 ;
        RECT 4.400 468.840 587.080 470.240 ;
        RECT 4.000 463.440 589.195 468.840 ;
        RECT 4.400 462.040 587.080 463.440 ;
        RECT 4.000 456.640 589.195 462.040 ;
        RECT 4.400 455.240 587.080 456.640 ;
        RECT 4.000 449.840 589.195 455.240 ;
        RECT 4.400 448.440 587.080 449.840 ;
        RECT 4.000 443.040 589.195 448.440 ;
        RECT 4.400 441.640 587.080 443.040 ;
        RECT 4.000 436.240 589.195 441.640 ;
        RECT 4.400 434.840 587.080 436.240 ;
        RECT 4.000 429.440 589.195 434.840 ;
        RECT 4.400 428.040 587.080 429.440 ;
        RECT 4.000 422.640 589.195 428.040 ;
        RECT 4.400 421.240 587.080 422.640 ;
        RECT 4.000 415.840 589.195 421.240 ;
        RECT 4.400 414.440 587.080 415.840 ;
        RECT 4.000 409.040 589.195 414.440 ;
        RECT 4.400 407.640 587.080 409.040 ;
        RECT 4.000 402.240 589.195 407.640 ;
        RECT 4.400 400.840 587.080 402.240 ;
        RECT 4.000 395.440 589.195 400.840 ;
        RECT 4.400 394.040 587.080 395.440 ;
        RECT 4.000 388.640 589.195 394.040 ;
        RECT 4.400 387.240 587.080 388.640 ;
        RECT 4.000 381.840 589.195 387.240 ;
        RECT 4.400 380.440 587.080 381.840 ;
        RECT 4.000 375.040 589.195 380.440 ;
        RECT 4.400 373.640 587.080 375.040 ;
        RECT 4.000 368.240 589.195 373.640 ;
        RECT 4.400 366.840 587.080 368.240 ;
        RECT 4.000 361.440 589.195 366.840 ;
        RECT 4.400 360.040 587.080 361.440 ;
        RECT 4.000 354.640 589.195 360.040 ;
        RECT 4.400 353.240 587.080 354.640 ;
        RECT 4.000 347.840 589.195 353.240 ;
        RECT 4.400 346.440 587.080 347.840 ;
        RECT 4.000 341.040 589.195 346.440 ;
        RECT 4.400 339.640 587.080 341.040 ;
        RECT 4.000 334.240 589.195 339.640 ;
        RECT 4.400 332.840 587.080 334.240 ;
        RECT 4.000 327.440 589.195 332.840 ;
        RECT 4.400 326.040 587.080 327.440 ;
        RECT 4.000 320.640 589.195 326.040 ;
        RECT 4.400 319.240 587.080 320.640 ;
        RECT 4.000 313.840 589.195 319.240 ;
        RECT 4.400 312.440 587.080 313.840 ;
        RECT 4.000 307.040 589.195 312.440 ;
        RECT 4.400 305.640 587.080 307.040 ;
        RECT 4.000 300.240 589.195 305.640 ;
        RECT 4.400 298.840 587.080 300.240 ;
        RECT 4.000 293.440 589.195 298.840 ;
        RECT 4.400 292.040 587.080 293.440 ;
        RECT 4.000 286.640 589.195 292.040 ;
        RECT 4.400 285.240 587.080 286.640 ;
        RECT 4.000 279.840 589.195 285.240 ;
        RECT 4.400 278.440 587.080 279.840 ;
        RECT 4.000 273.040 589.195 278.440 ;
        RECT 4.400 271.640 587.080 273.040 ;
        RECT 4.000 266.240 589.195 271.640 ;
        RECT 4.400 264.840 587.080 266.240 ;
        RECT 4.000 259.440 589.195 264.840 ;
        RECT 4.400 258.040 587.080 259.440 ;
        RECT 4.000 252.640 589.195 258.040 ;
        RECT 4.400 251.240 587.080 252.640 ;
        RECT 4.000 245.840 589.195 251.240 ;
        RECT 4.400 244.440 587.080 245.840 ;
        RECT 4.000 239.040 589.195 244.440 ;
        RECT 4.400 237.640 587.080 239.040 ;
        RECT 4.000 232.240 589.195 237.640 ;
        RECT 4.400 230.840 587.080 232.240 ;
        RECT 4.000 225.440 589.195 230.840 ;
        RECT 4.400 224.040 587.080 225.440 ;
        RECT 4.000 218.640 589.195 224.040 ;
        RECT 4.400 217.240 587.080 218.640 ;
        RECT 4.000 211.840 589.195 217.240 ;
        RECT 4.400 210.440 587.080 211.840 ;
        RECT 4.000 205.040 589.195 210.440 ;
        RECT 4.400 203.640 587.080 205.040 ;
        RECT 4.000 198.240 589.195 203.640 ;
        RECT 4.400 196.840 587.080 198.240 ;
        RECT 4.000 191.440 589.195 196.840 ;
        RECT 4.400 190.040 587.080 191.440 ;
        RECT 4.000 184.640 589.195 190.040 ;
        RECT 4.400 183.240 587.080 184.640 ;
        RECT 4.000 177.840 589.195 183.240 ;
        RECT 4.400 176.440 587.080 177.840 ;
        RECT 4.000 171.040 589.195 176.440 ;
        RECT 4.400 169.640 587.080 171.040 ;
        RECT 4.000 164.240 589.195 169.640 ;
        RECT 4.400 162.840 587.080 164.240 ;
        RECT 4.000 157.440 589.195 162.840 ;
        RECT 4.400 156.040 587.080 157.440 ;
        RECT 4.000 150.640 589.195 156.040 ;
        RECT 4.400 149.240 587.080 150.640 ;
        RECT 4.000 143.840 589.195 149.240 ;
        RECT 4.400 142.440 587.080 143.840 ;
        RECT 4.000 137.040 589.195 142.440 ;
        RECT 4.400 135.640 587.080 137.040 ;
        RECT 4.000 130.240 589.195 135.640 ;
        RECT 4.400 128.840 587.080 130.240 ;
        RECT 4.000 123.440 589.195 128.840 ;
        RECT 4.400 122.040 587.080 123.440 ;
        RECT 4.000 116.640 589.195 122.040 ;
        RECT 4.400 115.240 587.080 116.640 ;
        RECT 4.000 109.840 589.195 115.240 ;
        RECT 4.400 108.440 587.080 109.840 ;
        RECT 4.000 103.040 589.195 108.440 ;
        RECT 4.400 101.640 587.080 103.040 ;
        RECT 4.000 96.240 589.195 101.640 ;
        RECT 4.400 94.840 587.080 96.240 ;
        RECT 4.000 89.440 589.195 94.840 ;
        RECT 4.400 88.040 587.080 89.440 ;
        RECT 4.000 82.640 589.195 88.040 ;
        RECT 4.400 81.240 587.080 82.640 ;
        RECT 4.000 75.840 589.195 81.240 ;
        RECT 4.400 74.440 587.080 75.840 ;
        RECT 4.000 69.040 589.195 74.440 ;
        RECT 4.400 67.640 587.080 69.040 ;
        RECT 4.000 62.240 589.195 67.640 ;
        RECT 4.400 60.840 587.080 62.240 ;
        RECT 4.000 55.440 589.195 60.840 ;
        RECT 4.400 54.040 587.080 55.440 ;
        RECT 4.000 48.640 589.195 54.040 ;
        RECT 4.400 47.240 587.080 48.640 ;
        RECT 4.000 41.840 589.195 47.240 ;
        RECT 4.400 40.440 587.080 41.840 ;
        RECT 4.000 35.040 589.195 40.440 ;
        RECT 4.400 33.640 587.080 35.040 ;
        RECT 4.000 28.240 589.195 33.640 ;
        RECT 4.400 26.840 587.080 28.240 ;
        RECT 4.000 21.440 589.195 26.840 ;
        RECT 4.400 20.040 587.080 21.440 ;
        RECT 4.000 14.640 589.195 20.040 ;
        RECT 4.400 13.240 587.080 14.640 ;
        RECT 4.000 7.840 589.195 13.240 ;
        RECT 4.400 6.440 587.080 7.840 ;
        RECT 4.000 1.040 589.195 6.440 ;
        RECT 4.000 0.175 587.080 1.040 ;
      LAYER met4 ;
        RECT 9.495 590.880 579.305 600.945 ;
        RECT 9.495 10.240 20.640 590.880 ;
        RECT 23.040 10.240 97.440 590.880 ;
        RECT 99.840 10.240 174.240 590.880 ;
        RECT 176.640 10.240 251.040 590.880 ;
        RECT 253.440 10.240 327.840 590.880 ;
        RECT 330.240 10.240 404.640 590.880 ;
        RECT 407.040 10.240 481.440 590.880 ;
        RECT 483.840 10.240 558.240 590.880 ;
        RECT 560.640 10.240 579.305 590.880 ;
        RECT 9.495 5.615 579.305 10.240 ;
  END
END rvj1_caravel_soc
END LIBRARY

